magic
tech scmos
timestamp 1681696376
<< metal1 >>
rect -10 9 10 10
rect 9 -10 10 9
<< m2contact >>
rect -10 -10 9 9
<< metal2 >>
rect -10 9 10 10
rect 9 -10 10 9
<< end >>
