magic
tech scmos
timestamp 1683038052
<< metal1 >>
rect 14 1707 1750 1727
rect 38 1683 1726 1703
rect 14 1667 1750 1673
rect 506 1633 516 1636
rect 818 1633 828 1636
rect 418 1623 436 1626
rect 836 1623 853 1626
rect 908 1623 933 1626
rect 426 1616 429 1623
rect 132 1613 149 1616
rect 188 1613 205 1616
rect 412 1613 429 1616
rect 530 1613 540 1616
rect 914 1613 948 1616
rect 1212 1613 1228 1616
rect 1346 1613 1396 1616
rect 1540 1613 1557 1616
rect 1346 1607 1349 1613
rect 556 1603 573 1606
rect 770 1603 796 1606
rect 842 1603 860 1606
rect 884 1603 892 1606
rect 906 1603 940 1606
rect 1194 1603 1204 1606
rect 1354 1603 1388 1606
rect 1500 1603 1525 1606
rect 38 1567 1726 1573
rect 154 1533 164 1536
rect 212 1533 220 1536
rect 234 1533 244 1536
rect 282 1533 300 1536
rect 362 1533 380 1536
rect 778 1533 796 1536
rect 844 1533 861 1536
rect 906 1533 924 1536
rect 948 1533 1004 1536
rect 1018 1533 1068 1536
rect 1396 1533 1413 1536
rect 1426 1533 1436 1536
rect 1490 1533 1500 1536
rect 562 1526 565 1533
rect 1602 1526 1605 1533
rect 146 1523 172 1526
rect 186 1523 204 1526
rect 210 1523 228 1526
rect 284 1523 308 1526
rect 404 1523 429 1526
rect 468 1523 476 1526
rect 546 1523 556 1526
rect 562 1523 572 1526
rect 772 1523 789 1526
rect 804 1523 821 1526
rect 866 1523 876 1526
rect 890 1523 932 1526
rect 1002 1523 1012 1526
rect 1076 1523 1109 1526
rect 1402 1523 1428 1526
rect 1460 1523 1485 1526
rect 1508 1523 1525 1526
rect 1602 1523 1637 1526
rect 92 1513 101 1516
rect 850 1513 868 1516
rect 1562 1513 1580 1516
rect 90 1503 108 1506
rect 14 1467 1750 1473
rect 596 1433 613 1436
rect 778 1433 820 1436
rect 194 1423 204 1426
rect 562 1423 588 1426
rect 786 1423 804 1426
rect 828 1423 853 1426
rect 900 1423 933 1426
rect 1138 1423 1156 1426
rect 74 1413 133 1416
rect 210 1413 236 1416
rect 266 1413 292 1416
rect 338 1413 348 1416
rect 378 1413 404 1416
rect 442 1413 452 1416
rect 458 1413 493 1416
rect 500 1413 509 1416
rect 732 1413 741 1416
rect 338 1407 341 1413
rect 116 1403 141 1406
rect 538 1403 548 1406
rect 618 1403 628 1406
rect 538 1395 541 1403
rect 738 1395 741 1413
rect 754 1403 757 1414
rect 762 1407 765 1416
rect 772 1413 797 1416
rect 860 1413 884 1416
rect 970 1413 996 1416
rect 1002 1413 1020 1416
rect 1420 1413 1445 1416
rect 1452 1413 1485 1416
rect 1684 1413 1693 1416
rect 1442 1407 1445 1413
rect 834 1403 852 1406
rect 906 1403 932 1406
rect 962 1403 988 1406
rect 1124 1403 1149 1406
rect 1186 1403 1260 1406
rect 1428 1403 1437 1406
rect 38 1367 1726 1373
rect 898 1336 901 1346
rect 170 1333 196 1336
rect 298 1333 308 1336
rect 340 1333 348 1336
rect 540 1333 557 1336
rect 754 1333 764 1336
rect 882 1333 916 1336
rect 954 1333 964 1336
rect 1194 1333 1212 1336
rect 1322 1333 1349 1336
rect 1386 1333 1420 1336
rect 130 1326 133 1333
rect 130 1323 140 1326
rect 178 1323 204 1326
rect 226 1323 229 1333
rect 282 1326 285 1333
rect 394 1326 397 1333
rect 754 1326 757 1333
rect 268 1323 285 1326
rect 298 1323 316 1326
rect 356 1323 397 1326
rect 418 1323 436 1326
rect 554 1323 564 1326
rect 748 1323 757 1326
rect 772 1323 781 1326
rect 788 1323 821 1326
rect 868 1323 877 1326
rect 882 1323 885 1333
rect 940 1323 965 1326
rect 1130 1323 1156 1326
rect 1258 1323 1284 1326
rect 1346 1325 1349 1333
rect 1380 1323 1413 1326
rect 1538 1323 1548 1326
rect 1620 1323 1636 1326
rect 298 1315 301 1323
rect 418 1315 421 1323
rect 796 1313 860 1316
rect 1578 1313 1604 1316
rect 14 1267 1750 1273
rect 514 1233 524 1236
rect 66 1213 84 1216
rect 220 1213 229 1216
rect 268 1213 285 1216
rect 346 1213 356 1216
rect 418 1213 436 1216
rect 538 1213 548 1216
rect 612 1213 629 1216
rect 796 1213 805 1216
rect 874 1213 917 1216
rect 948 1213 981 1216
rect 1116 1213 1125 1216
rect 1140 1213 1164 1216
rect 1218 1213 1228 1216
rect 1258 1213 1269 1216
rect 1292 1213 1301 1216
rect 1314 1213 1324 1216
rect 1418 1213 1445 1216
rect 1532 1213 1541 1216
rect 1684 1213 1693 1216
rect 226 1207 229 1213
rect 874 1207 877 1213
rect 914 1206 917 1213
rect 1258 1207 1261 1213
rect 1314 1207 1317 1213
rect 1442 1207 1445 1213
rect 90 1203 100 1206
rect 482 1203 492 1206
rect 564 1203 597 1206
rect 820 1203 828 1206
rect 914 1203 932 1206
rect 962 1203 980 1206
rect 1098 1203 1108 1206
rect 1202 1203 1220 1206
rect 1354 1203 1364 1206
rect 38 1167 1726 1173
rect 84 1133 93 1136
rect 194 1126 197 1135
rect 810 1133 820 1136
rect 842 1133 852 1136
rect 1058 1133 1084 1136
rect 1322 1133 1332 1136
rect 1386 1133 1428 1136
rect 1450 1133 1508 1136
rect 1660 1133 1693 1136
rect 66 1123 76 1126
rect 188 1123 197 1126
rect 354 1123 380 1126
rect 410 1123 436 1126
rect 732 1123 797 1126
rect 802 1123 812 1126
rect 844 1123 853 1126
rect 884 1123 900 1126
rect 954 1123 980 1126
rect 1060 1123 1085 1126
rect 1228 1123 1253 1126
rect 1324 1123 1333 1126
rect 1410 1123 1420 1126
rect 1452 1123 1477 1126
rect 1612 1123 1621 1126
rect 1636 1123 1652 1126
rect 674 1113 716 1116
rect 14 1067 1750 1073
rect 1618 1033 1637 1036
rect 90 1013 100 1016
rect 482 1013 492 1016
rect 82 1003 108 1006
rect 124 1003 133 1006
rect 252 1003 285 1006
rect 308 1003 324 1006
rect 460 1003 493 1006
rect 522 1003 525 1014
rect 540 1013 556 1016
rect 578 1013 660 1016
rect 794 1013 804 1016
rect 844 1013 861 1016
rect 900 1013 909 1016
rect 986 1006 989 1014
rect 1020 1013 1045 1016
rect 1218 1013 1236 1016
rect 1348 1013 1357 1016
rect 1474 1013 1500 1016
rect 1572 1013 1580 1016
rect 1676 1013 1765 1016
rect 572 1003 637 1006
rect 642 1003 668 1006
rect 940 1003 949 1006
rect 972 1003 989 1006
rect 1012 1003 1021 1006
rect 1026 1003 1044 1006
rect 1154 1003 1164 1006
rect 1212 1003 1229 1006
rect 1306 1003 1324 1006
rect 1346 1003 1364 1006
rect 1498 1003 1508 1006
rect 1524 1003 1541 1006
rect 1578 1003 1588 1006
rect 1618 1003 1652 1006
rect 38 967 1726 973
rect 1146 936 1149 946
rect 1202 943 1228 946
rect 82 933 116 936
rect 284 933 293 936
rect 460 933 485 936
rect 514 933 572 936
rect 1012 933 1021 936
rect 1138 933 1172 936
rect 1218 933 1236 936
rect 1242 933 1276 936
rect 1298 933 1356 936
rect 1378 933 1412 936
rect 1458 933 1532 936
rect 1548 933 1589 936
rect 1612 933 1629 936
rect 1642 933 1660 936
rect 314 926 317 933
rect 66 923 108 926
rect 140 923 157 926
rect 228 923 269 926
rect 282 923 308 926
rect 314 923 333 926
rect 346 923 349 933
rect 466 923 484 926
rect 516 923 533 926
rect 546 923 580 926
rect 690 923 700 926
rect 884 923 901 926
rect 980 923 989 926
rect 1060 923 1101 926
rect 1138 925 1141 933
rect 1146 923 1164 926
rect 1250 923 1268 926
rect 1300 923 1349 926
rect 1354 923 1364 926
rect 1420 923 1436 926
rect 1490 923 1524 926
rect 1650 923 1668 926
rect 1684 923 1693 926
rect 146 913 212 916
rect 1452 913 1477 916
rect 14 867 1750 873
rect 1148 823 1157 826
rect 1154 816 1157 823
rect 1282 816 1285 826
rect 66 813 76 816
rect 108 813 116 816
rect 402 803 405 814
rect 410 807 413 816
rect 540 813 549 816
rect 666 803 669 814
rect 682 813 700 816
rect 706 813 716 816
rect 860 813 885 816
rect 1154 813 1172 816
rect 1196 813 1205 816
rect 1218 813 1244 816
rect 1282 813 1293 816
rect 1340 813 1357 816
rect 1434 813 1460 816
rect 1612 813 1629 816
rect 1290 807 1293 813
rect 1674 807 1677 816
rect 1684 813 1693 816
rect 676 803 692 806
rect 1082 803 1100 806
rect 1194 803 1204 806
rect 1260 803 1285 806
rect 1420 803 1461 806
rect 1484 803 1509 806
rect 1514 803 1532 806
rect 1548 803 1581 806
rect 1618 803 1660 806
rect 1690 803 1693 813
rect 1218 793 1244 796
rect 38 767 1726 773
rect 596 743 605 746
rect 538 733 564 736
rect 570 733 588 736
rect 628 733 637 736
rect 642 733 676 736
rect 274 726 277 733
rect 282 726 285 733
rect 66 723 76 726
rect 204 723 213 726
rect 274 723 285 726
rect 530 723 533 733
rect 682 726 685 744
rect 738 733 748 736
rect 572 723 580 726
rect 594 723 620 726
rect 682 723 700 726
rect 706 723 709 733
rect 714 723 724 726
rect 730 723 733 733
rect 754 726 757 744
rect 1210 743 1260 746
rect 762 733 772 736
rect 810 733 836 736
rect 930 733 940 736
rect 1196 733 1229 736
rect 1274 733 1285 736
rect 1314 733 1348 736
rect 1530 733 1557 736
rect 1594 733 1604 736
rect 906 726 909 733
rect 754 723 772 726
rect 906 723 917 726
rect 978 723 996 726
rect 1010 723 1044 726
rect 1138 723 1156 726
rect 1204 723 1221 726
rect 1282 725 1285 733
rect 1316 723 1325 726
rect 1330 723 1340 726
rect 1434 723 1460 726
rect 1530 725 1533 733
rect 1538 723 1556 726
rect 14 667 1750 673
rect 1548 623 1557 626
rect 1604 623 1613 626
rect 66 613 108 616
rect 146 613 180 616
rect 212 613 221 616
rect 338 613 356 616
rect 500 613 509 616
rect 572 613 581 616
rect 634 613 652 616
rect 794 613 812 616
rect 940 613 957 616
rect 996 613 1012 616
rect 1044 613 1053 616
rect 1074 613 1084 616
rect 1212 613 1228 616
rect 1356 613 1380 616
rect 1394 613 1404 616
rect 1516 613 1532 616
rect 1546 613 1565 616
rect 1572 613 1588 616
rect 1562 607 1565 613
rect 82 603 116 606
rect 332 603 357 606
rect 524 603 564 606
rect 570 603 588 606
rect 612 603 637 606
rect 642 603 652 606
rect 706 603 732 606
rect 770 603 812 606
rect 874 603 908 606
rect 946 603 964 606
rect 1178 603 1204 606
rect 1604 603 1629 606
rect 538 593 556 596
rect 708 593 717 596
rect 874 593 877 603
rect 38 567 1726 573
rect 298 533 308 536
rect 546 533 556 536
rect 618 533 652 536
rect 690 533 708 536
rect 746 533 756 536
rect 794 533 804 536
rect 842 533 852 536
rect 922 533 932 536
rect 986 533 996 536
rect 546 526 549 533
rect 66 523 108 526
rect 140 523 157 526
rect 220 523 301 526
rect 532 523 549 526
rect 564 523 573 526
rect 634 523 652 526
rect 684 523 693 526
rect 698 523 708 526
rect 842 523 852 526
rect 924 523 948 526
rect 978 523 981 533
rect 1028 523 1036 526
rect 1132 523 1141 526
rect 1188 523 1197 526
rect 1340 523 1357 526
rect 1436 523 1445 526
rect 1684 523 1701 526
rect 146 513 204 516
rect 14 467 1750 473
rect 66 413 84 416
rect 322 413 332 416
rect 394 406 397 414
rect 402 413 476 416
rect 546 413 556 416
rect 602 413 628 416
rect 700 413 741 416
rect 762 413 796 416
rect 876 413 885 416
rect 340 403 365 406
rect 394 403 421 406
rect 484 403 541 406
rect 546 393 549 413
rect 588 403 621 406
rect 700 403 709 406
rect 738 395 741 413
rect 748 403 797 406
rect 804 403 852 406
rect 898 405 901 416
rect 948 413 981 416
rect 1012 413 1021 416
rect 1066 413 1092 416
rect 1124 413 1133 416
rect 1170 413 1204 416
rect 1324 413 1333 416
rect 1354 413 1364 416
rect 1556 413 1573 416
rect 1684 413 1693 416
rect 978 406 981 413
rect 932 403 940 406
rect 978 403 996 406
rect 1074 403 1100 406
rect 1122 403 1132 406
rect 1338 403 1356 406
rect 1410 403 1436 406
rect 1570 403 1580 406
rect 954 393 988 396
rect 1410 393 1413 403
rect 1570 383 1573 403
rect 38 367 1726 373
rect 116 333 133 336
rect 588 333 605 336
rect 684 333 701 336
rect 740 333 757 336
rect 796 333 837 336
rect 844 333 853 336
rect 850 326 853 333
rect 874 326 877 344
rect 82 323 92 326
rect 164 323 173 326
rect 188 323 204 326
rect 620 323 645 326
rect 754 323 764 326
rect 802 323 836 326
rect 850 323 861 326
rect 868 323 877 326
rect 890 325 893 336
rect 1154 333 1172 336
rect 1242 333 1252 336
rect 1274 333 1332 336
rect 1370 333 1404 336
rect 1684 333 1693 336
rect 1554 326 1557 333
rect 898 323 908 326
rect 1028 323 1044 326
rect 1212 323 1229 326
rect 1260 323 1269 326
rect 1290 323 1324 326
rect 1356 323 1381 326
rect 1540 323 1557 326
rect 14 267 1750 273
rect 66 213 84 216
rect 212 213 228 216
rect 348 213 364 216
rect 452 213 484 216
rect 580 213 589 216
rect 628 213 637 216
rect 812 213 845 216
rect 964 213 1004 216
rect 1170 213 1180 216
rect 410 203 428 206
rect 450 203 460 206
rect 508 203 516 206
rect 580 203 589 206
rect 628 203 637 206
rect 676 203 693 206
rect 732 203 749 206
rect 788 203 797 206
rect 866 195 869 206
rect 884 203 901 206
rect 908 203 956 206
rect 970 203 996 206
rect 1530 203 1533 214
rect 1562 203 1565 214
rect 1684 203 1693 206
rect 38 167 1726 173
rect 364 143 397 146
rect 394 136 397 143
rect 786 136 789 146
rect 316 133 333 136
rect 356 133 389 136
rect 394 133 404 136
rect 500 133 509 136
rect 668 133 685 136
rect 748 133 804 136
rect 450 126 453 133
rect 866 126 869 144
rect 876 133 893 136
rect 900 133 933 136
rect 1052 133 1061 136
rect 1586 133 1596 136
rect 290 123 308 126
rect 394 123 420 126
rect 450 123 492 126
rect 522 123 540 126
rect 586 123 596 126
rect 628 123 636 126
rect 674 123 692 126
rect 724 123 741 126
rect 828 123 869 126
rect 884 123 892 126
rect 1458 123 1468 126
rect 1604 123 1685 126
rect 14 67 1750 73
rect 38 37 1726 57
rect 14 13 1750 33
<< metal2 >>
rect 14 13 34 1727
rect 38 37 58 1703
rect 74 1533 85 1536
rect 106 1533 109 1606
rect 114 1533 125 1536
rect 146 1533 149 1616
rect 202 1573 205 1616
rect 82 1506 85 1526
rect 98 1523 109 1526
rect 82 1503 93 1506
rect 98 1486 101 1516
rect 90 1483 101 1486
rect 74 1226 77 1416
rect 90 1336 93 1483
rect 106 1406 109 1523
rect 114 1513 117 1533
rect 122 1456 125 1526
rect 130 1513 133 1526
rect 138 1523 149 1526
rect 82 1333 93 1336
rect 98 1403 109 1406
rect 118 1453 125 1456
rect 118 1406 121 1453
rect 130 1413 133 1446
rect 118 1403 125 1406
rect 90 1236 93 1326
rect 98 1303 101 1403
rect 122 1386 125 1403
rect 138 1393 141 1523
rect 146 1423 149 1516
rect 154 1503 157 1536
rect 210 1533 213 1616
rect 234 1533 237 1576
rect 250 1543 261 1546
rect 178 1503 181 1516
rect 186 1513 189 1526
rect 154 1433 157 1446
rect 162 1413 165 1426
rect 122 1383 141 1386
rect 106 1333 125 1336
rect 114 1313 117 1326
rect 90 1233 101 1236
rect 74 1223 93 1226
rect 66 1123 69 1216
rect 74 1203 93 1206
rect 98 1196 101 1233
rect 90 1193 101 1196
rect 106 1193 109 1216
rect 122 1213 125 1333
rect 130 1303 133 1316
rect 90 1143 93 1193
rect 90 1113 93 1136
rect 106 1133 109 1146
rect 130 1113 133 1126
rect 138 1083 141 1383
rect 146 1333 149 1346
rect 162 1343 165 1396
rect 170 1333 173 1426
rect 178 1343 181 1426
rect 186 1423 189 1436
rect 194 1423 197 1516
rect 210 1503 213 1526
rect 250 1506 253 1543
rect 266 1536 269 1616
rect 290 1593 293 1606
rect 258 1533 269 1536
rect 258 1523 261 1533
rect 234 1503 253 1506
rect 274 1503 277 1536
rect 162 1213 165 1326
rect 178 1323 181 1336
rect 186 1313 189 1336
rect 194 1333 197 1416
rect 202 1413 213 1416
rect 234 1376 237 1503
rect 282 1486 285 1576
rect 278 1483 285 1486
rect 266 1376 269 1416
rect 234 1373 253 1376
rect 250 1353 253 1373
rect 258 1373 269 1376
rect 226 1306 229 1326
rect 218 1303 229 1306
rect 234 1303 237 1326
rect 218 1246 221 1303
rect 218 1243 229 1246
rect 226 1213 229 1243
rect 242 1216 245 1336
rect 250 1323 253 1336
rect 258 1333 261 1373
rect 278 1366 281 1483
rect 278 1363 285 1366
rect 274 1333 277 1346
rect 250 1223 253 1236
rect 194 1133 197 1166
rect 202 1123 205 1186
rect 234 1163 237 1216
rect 242 1213 253 1216
rect 250 1173 253 1213
rect 258 1203 261 1226
rect 266 1183 269 1326
rect 282 1243 285 1363
rect 290 1313 293 1526
rect 306 1513 309 1526
rect 298 1333 301 1346
rect 290 1236 293 1296
rect 274 1233 293 1236
rect 274 1223 277 1233
rect 282 1213 285 1226
rect 290 1213 293 1233
rect 298 1206 301 1316
rect 306 1293 309 1356
rect 314 1243 317 1596
rect 330 1593 333 1636
rect 322 1533 325 1586
rect 354 1583 357 1616
rect 362 1536 365 1546
rect 346 1533 365 1536
rect 322 1503 325 1516
rect 330 1513 333 1526
rect 338 1513 341 1526
rect 346 1503 349 1533
rect 354 1503 357 1516
rect 322 1333 325 1386
rect 330 1323 333 1436
rect 338 1413 341 1426
rect 378 1423 381 1566
rect 418 1553 421 1740
rect 466 1636 469 1646
rect 450 1633 469 1636
rect 442 1576 445 1616
rect 458 1613 461 1626
rect 434 1573 445 1576
rect 426 1533 429 1566
rect 426 1493 429 1526
rect 434 1496 437 1573
rect 442 1533 445 1546
rect 450 1503 453 1596
rect 434 1493 445 1496
rect 378 1383 381 1416
rect 442 1413 445 1493
rect 450 1406 453 1426
rect 458 1413 461 1606
rect 466 1536 469 1633
rect 482 1633 501 1636
rect 506 1633 509 1646
rect 530 1633 533 1740
rect 730 1656 733 1740
rect 722 1653 733 1656
rect 474 1583 477 1616
rect 482 1603 485 1633
rect 490 1613 493 1626
rect 498 1623 501 1633
rect 506 1613 509 1626
rect 522 1613 525 1626
rect 530 1613 533 1626
rect 490 1603 501 1606
rect 530 1593 533 1606
rect 466 1533 485 1536
rect 490 1513 493 1526
rect 498 1523 501 1536
rect 498 1513 517 1516
rect 466 1406 469 1496
rect 426 1383 429 1406
rect 442 1403 453 1406
rect 458 1403 469 1406
rect 490 1403 493 1416
rect 338 1323 341 1336
rect 354 1323 357 1346
rect 306 1216 309 1226
rect 314 1223 317 1236
rect 306 1213 317 1216
rect 322 1213 325 1316
rect 394 1303 397 1326
rect 402 1283 405 1326
rect 282 1203 301 1206
rect 306 1153 309 1206
rect 314 1183 317 1213
rect 330 1163 333 1236
rect 338 1213 341 1226
rect 346 1213 349 1226
rect 346 1183 349 1206
rect 210 1133 229 1136
rect 218 1113 221 1126
rect 226 1123 229 1133
rect 282 1123 285 1146
rect 306 1123 309 1136
rect 322 1133 325 1146
rect 330 1126 333 1156
rect 346 1133 349 1176
rect 322 1123 333 1126
rect 322 1113 325 1123
rect 66 913 69 926
rect 66 813 69 826
rect 82 786 85 1006
rect 90 993 93 1016
rect 114 1013 117 1046
rect 130 1013 133 1026
rect 98 896 101 926
rect 122 916 125 926
rect 130 923 133 1006
rect 146 956 149 1016
rect 162 1013 165 1036
rect 202 1013 205 1026
rect 226 966 229 1066
rect 242 1013 245 1026
rect 222 963 229 966
rect 146 953 157 956
rect 122 913 149 916
rect 154 903 157 953
rect 98 893 109 896
rect 106 836 109 893
rect 90 813 93 836
rect 98 833 109 836
rect 78 783 85 786
rect 66 673 69 726
rect 78 626 81 783
rect 98 766 101 833
rect 106 793 109 816
rect 170 803 173 816
rect 90 763 101 766
rect 66 613 69 626
rect 78 623 85 626
rect 82 603 85 623
rect 90 593 93 763
rect 106 613 109 676
rect 122 613 125 636
rect 130 626 133 726
rect 154 636 157 746
rect 178 733 181 776
rect 194 743 197 856
rect 210 843 213 936
rect 222 876 225 963
rect 222 873 229 876
rect 226 853 229 873
rect 210 823 213 836
rect 210 723 213 806
rect 218 646 221 766
rect 226 753 229 816
rect 234 763 237 956
rect 250 736 253 1086
rect 338 1046 341 1126
rect 330 1043 341 1046
rect 282 993 285 1006
rect 266 916 269 926
rect 274 923 277 976
rect 290 933 293 1016
rect 322 1003 325 1026
rect 330 996 333 1043
rect 354 1023 357 1166
rect 362 1123 365 1246
rect 370 1213 373 1226
rect 378 1213 381 1246
rect 418 1213 421 1336
rect 426 1303 429 1316
rect 442 1243 445 1403
rect 498 1336 501 1513
rect 522 1506 525 1536
rect 506 1503 525 1506
rect 530 1493 533 1586
rect 538 1526 541 1616
rect 554 1613 557 1626
rect 570 1603 573 1626
rect 586 1603 589 1616
rect 610 1613 613 1626
rect 546 1533 557 1536
rect 538 1523 549 1526
rect 546 1503 549 1516
rect 554 1446 557 1533
rect 562 1513 565 1526
rect 626 1496 629 1546
rect 666 1543 669 1616
rect 682 1536 685 1616
rect 706 1603 709 1616
rect 722 1566 725 1653
rect 818 1626 821 1636
rect 722 1563 733 1566
rect 650 1523 653 1536
rect 666 1523 669 1536
rect 674 1533 685 1536
rect 626 1493 637 1496
rect 546 1443 557 1446
rect 506 1423 525 1426
rect 506 1413 509 1423
rect 490 1333 501 1336
rect 498 1286 501 1326
rect 506 1296 509 1406
rect 514 1403 517 1416
rect 522 1346 525 1423
rect 522 1343 533 1346
rect 514 1323 517 1336
rect 522 1313 525 1336
rect 530 1323 533 1343
rect 538 1316 541 1416
rect 546 1403 549 1443
rect 562 1423 565 1456
rect 554 1333 557 1416
rect 602 1413 605 1446
rect 610 1433 621 1436
rect 594 1346 597 1366
rect 594 1343 601 1346
rect 538 1313 549 1316
rect 514 1296 517 1306
rect 506 1293 517 1296
rect 498 1283 509 1286
rect 498 1213 501 1226
rect 506 1223 509 1283
rect 514 1233 517 1293
rect 514 1213 517 1226
rect 530 1213 533 1226
rect 538 1213 541 1226
rect 546 1206 549 1313
rect 554 1303 557 1326
rect 598 1286 601 1343
rect 594 1283 601 1286
rect 562 1213 565 1226
rect 370 1133 373 1206
rect 458 1176 461 1206
rect 434 1173 461 1176
rect 434 1156 437 1173
rect 426 1153 437 1156
rect 410 1123 413 1136
rect 426 1096 429 1153
rect 458 1123 461 1166
rect 482 1123 485 1206
rect 538 1203 549 1206
rect 570 1186 573 1226
rect 594 1203 597 1283
rect 562 1183 573 1186
rect 426 1093 437 1096
rect 314 993 333 996
rect 330 933 333 993
rect 346 963 349 1016
rect 354 1013 365 1016
rect 410 1013 413 1026
rect 434 1003 437 1093
rect 450 1013 453 1026
rect 474 966 477 1016
rect 482 1003 485 1016
rect 490 996 493 1006
rect 498 1003 501 1016
rect 490 993 501 996
rect 506 993 509 1016
rect 474 963 493 966
rect 450 926 453 946
rect 282 916 285 926
rect 266 913 285 916
rect 330 923 341 926
rect 274 813 277 846
rect 242 733 253 736
rect 242 686 245 733
rect 258 703 261 726
rect 266 723 269 756
rect 210 643 221 646
rect 234 683 245 686
rect 154 633 161 636
rect 130 623 149 626
rect 130 613 141 616
rect 146 613 149 623
rect 66 513 69 526
rect 114 516 117 606
rect 106 513 117 516
rect 122 516 125 526
rect 130 523 133 606
rect 158 576 161 633
rect 194 623 197 636
rect 186 603 189 616
rect 210 606 213 643
rect 218 613 221 626
rect 194 603 205 606
rect 210 603 221 606
rect 218 586 221 603
rect 218 583 229 586
rect 158 573 173 576
rect 122 513 149 516
rect 66 413 69 476
rect 106 466 109 513
rect 106 463 117 466
rect 114 446 117 463
rect 114 443 121 446
rect 118 376 121 443
rect 114 373 121 376
rect 98 333 101 356
rect 114 353 117 373
rect 130 333 133 506
rect 154 473 157 526
rect 170 446 173 573
rect 162 443 173 446
rect 138 413 141 436
rect 138 333 141 356
rect 154 333 157 346
rect 82 303 85 326
rect 106 293 109 326
rect 66 213 69 276
rect 82 123 85 226
rect 122 223 125 326
rect 130 313 133 326
rect 146 316 149 326
rect 162 323 165 443
rect 170 333 181 336
rect 170 323 181 326
rect 146 313 173 316
rect 138 213 141 226
rect 162 133 165 306
rect 178 273 181 323
rect 194 303 197 476
rect 202 423 205 536
rect 226 473 229 583
rect 234 566 237 683
rect 258 603 261 616
rect 274 603 277 776
rect 330 763 333 923
rect 346 903 349 926
rect 338 803 341 816
rect 346 803 349 826
rect 354 813 357 926
rect 362 813 365 926
rect 450 923 469 926
rect 354 753 357 796
rect 362 783 365 806
rect 370 746 373 816
rect 378 773 381 866
rect 386 813 389 826
rect 394 813 405 816
rect 410 813 413 906
rect 474 903 477 946
rect 482 913 485 936
rect 490 863 493 963
rect 498 923 501 993
rect 514 966 517 1006
rect 506 963 517 966
rect 506 933 509 963
rect 514 923 517 936
rect 522 843 525 1006
rect 530 943 533 1056
rect 530 836 533 926
rect 522 833 533 836
rect 522 816 525 833
rect 386 796 389 806
rect 394 803 397 813
rect 386 793 397 796
rect 370 743 389 746
rect 394 733 397 793
rect 402 773 405 806
rect 410 743 413 806
rect 418 793 421 816
rect 426 786 429 816
rect 514 813 525 816
rect 538 813 541 1136
rect 562 1063 565 1183
rect 602 1163 605 1246
rect 610 1133 613 1426
rect 618 1403 621 1433
rect 634 1413 637 1493
rect 618 1186 621 1396
rect 642 1226 645 1386
rect 650 1376 653 1516
rect 674 1513 677 1533
rect 650 1373 669 1376
rect 634 1223 645 1226
rect 626 1206 629 1216
rect 634 1213 637 1223
rect 626 1203 645 1206
rect 618 1183 625 1186
rect 622 1126 625 1183
rect 650 1173 653 1216
rect 658 1203 661 1216
rect 666 1196 669 1373
rect 674 1363 677 1416
rect 682 1383 685 1526
rect 698 1456 701 1546
rect 730 1543 733 1563
rect 722 1513 725 1526
rect 746 1523 749 1536
rect 762 1513 765 1626
rect 802 1623 813 1626
rect 818 1623 829 1626
rect 770 1536 773 1606
rect 770 1533 781 1536
rect 694 1453 701 1456
rect 694 1376 697 1453
rect 722 1413 733 1416
rect 746 1403 749 1426
rect 762 1416 765 1506
rect 778 1423 781 1436
rect 786 1423 789 1536
rect 802 1506 805 1623
rect 818 1566 821 1616
rect 826 1606 829 1623
rect 850 1613 853 1626
rect 858 1623 861 1740
rect 970 1726 973 1740
rect 962 1723 973 1726
rect 962 1656 965 1723
rect 962 1653 973 1656
rect 826 1603 833 1606
rect 810 1563 821 1566
rect 810 1513 813 1563
rect 830 1546 833 1603
rect 842 1593 845 1606
rect 818 1533 821 1546
rect 826 1543 833 1546
rect 818 1516 821 1526
rect 826 1523 829 1543
rect 818 1513 845 1516
rect 850 1513 853 1526
rect 802 1503 813 1506
rect 754 1413 765 1416
rect 694 1373 701 1376
rect 690 1313 693 1326
rect 698 1306 701 1373
rect 754 1333 757 1406
rect 778 1323 781 1346
rect 794 1313 797 1436
rect 802 1396 805 1426
rect 810 1416 813 1503
rect 850 1423 853 1446
rect 810 1413 837 1416
rect 858 1413 861 1536
rect 866 1523 869 1616
rect 882 1613 885 1626
rect 898 1593 901 1616
rect 906 1613 917 1616
rect 874 1533 885 1536
rect 866 1423 869 1436
rect 834 1403 837 1413
rect 802 1393 809 1396
rect 806 1306 809 1393
rect 874 1333 877 1526
rect 890 1513 893 1526
rect 898 1506 901 1546
rect 890 1503 901 1506
rect 906 1503 909 1606
rect 922 1546 925 1636
rect 970 1633 973 1653
rect 986 1626 989 1740
rect 930 1606 933 1626
rect 962 1616 965 1626
rect 954 1613 965 1616
rect 970 1623 989 1626
rect 930 1603 937 1606
rect 918 1543 925 1546
rect 890 1416 893 1503
rect 918 1496 921 1543
rect 934 1536 937 1603
rect 914 1493 921 1496
rect 930 1533 937 1536
rect 886 1413 893 1416
rect 886 1356 889 1413
rect 886 1353 893 1356
rect 890 1336 893 1353
rect 898 1343 901 1406
rect 906 1403 909 1416
rect 914 1336 917 1493
rect 930 1446 933 1533
rect 946 1513 949 1596
rect 954 1556 957 1613
rect 962 1573 965 1606
rect 954 1553 961 1556
rect 958 1506 961 1553
rect 954 1503 961 1506
rect 930 1443 941 1446
rect 954 1443 957 1503
rect 930 1423 933 1436
rect 938 1413 941 1443
rect 890 1333 901 1336
rect 658 1193 669 1196
rect 690 1303 701 1306
rect 802 1303 809 1306
rect 818 1306 821 1326
rect 874 1306 877 1326
rect 818 1303 829 1306
rect 578 1053 581 1126
rect 618 1123 625 1126
rect 618 1076 621 1123
rect 610 1073 621 1076
rect 570 1023 573 1046
rect 546 953 549 1016
rect 578 1013 581 1036
rect 610 996 613 1073
rect 634 1003 637 1126
rect 658 1083 661 1193
rect 674 1013 677 1116
rect 690 1013 693 1303
rect 802 1233 805 1303
rect 826 1246 829 1303
rect 818 1243 829 1246
rect 866 1303 877 1306
rect 866 1246 869 1303
rect 866 1243 877 1246
rect 714 1213 717 1226
rect 738 1143 741 1216
rect 754 1213 757 1226
rect 802 1213 805 1226
rect 714 1126 717 1136
rect 714 1123 725 1126
rect 610 993 621 996
rect 546 906 549 926
rect 586 913 589 926
rect 618 923 621 993
rect 642 963 645 1006
rect 674 943 677 1006
rect 682 973 685 1006
rect 706 1003 709 1086
rect 722 1066 725 1123
rect 722 1063 733 1066
rect 730 1013 733 1063
rect 738 1013 741 1136
rect 746 1116 749 1176
rect 754 1133 757 1196
rect 762 1146 765 1206
rect 770 1163 773 1206
rect 762 1143 773 1146
rect 746 1113 753 1116
rect 750 1026 753 1113
rect 746 1023 753 1026
rect 746 1003 749 1023
rect 770 963 773 1143
rect 786 1006 789 1016
rect 794 1013 797 1126
rect 802 1123 805 1186
rect 818 1153 821 1243
rect 842 1213 853 1216
rect 826 1173 829 1206
rect 874 1186 877 1243
rect 810 1036 813 1136
rect 802 1033 813 1036
rect 786 1003 797 1006
rect 690 936 693 956
rect 794 953 797 1003
rect 802 986 805 1033
rect 818 1003 821 1146
rect 826 1143 845 1146
rect 826 1123 829 1143
rect 834 1046 837 1136
rect 842 1133 845 1143
rect 850 1123 853 1186
rect 866 1183 877 1186
rect 858 1106 861 1126
rect 854 1103 861 1106
rect 834 1043 845 1046
rect 842 996 845 1043
rect 854 1036 857 1103
rect 854 1033 861 1036
rect 858 1013 861 1033
rect 866 1013 869 1183
rect 874 1113 877 1176
rect 882 1163 885 1326
rect 898 1246 901 1333
rect 910 1333 917 1336
rect 910 1286 913 1333
rect 922 1296 925 1326
rect 946 1316 949 1336
rect 954 1333 957 1416
rect 970 1413 973 1623
rect 978 1593 981 1606
rect 986 1533 989 1616
rect 994 1516 997 1616
rect 1090 1603 1093 1616
rect 986 1513 997 1516
rect 986 1416 989 1513
rect 986 1413 997 1416
rect 1002 1413 1005 1526
rect 1018 1446 1021 1596
rect 1082 1533 1085 1596
rect 1098 1593 1101 1616
rect 1106 1513 1109 1526
rect 1010 1443 1021 1446
rect 962 1333 965 1406
rect 994 1393 997 1413
rect 1010 1403 1013 1443
rect 1114 1436 1117 1526
rect 1122 1503 1125 1536
rect 1114 1433 1125 1436
rect 1122 1416 1125 1433
rect 946 1313 957 1316
rect 962 1313 965 1326
rect 922 1293 933 1296
rect 910 1283 917 1286
rect 894 1243 901 1246
rect 894 1196 897 1243
rect 894 1193 901 1196
rect 834 993 845 996
rect 802 983 821 986
rect 794 943 813 946
rect 682 913 685 936
rect 690 933 701 936
rect 546 903 557 906
rect 554 846 557 903
rect 546 843 557 846
rect 546 813 549 843
rect 514 793 517 813
rect 418 783 429 786
rect 522 783 525 806
rect 530 803 541 806
rect 402 733 413 736
rect 418 733 421 783
rect 426 743 429 776
rect 282 703 285 726
rect 290 713 293 726
rect 298 656 301 726
rect 394 706 397 726
rect 402 713 405 726
rect 498 723 501 746
rect 378 703 397 706
rect 298 653 305 656
rect 302 576 305 653
rect 314 633 333 636
rect 314 613 317 633
rect 322 613 325 626
rect 298 573 305 576
rect 234 563 245 566
rect 242 466 245 563
rect 298 533 301 573
rect 314 543 317 606
rect 330 603 333 633
rect 338 603 341 616
rect 362 613 373 616
rect 354 553 357 606
rect 362 593 365 606
rect 298 506 301 526
rect 378 523 381 703
rect 386 596 389 616
rect 394 603 397 666
rect 514 663 517 726
rect 522 723 525 746
rect 538 733 541 796
rect 530 703 533 726
rect 538 696 541 726
rect 530 693 541 696
rect 506 623 525 626
rect 386 593 405 596
rect 298 503 317 506
rect 226 463 245 466
rect 210 323 213 336
rect 178 213 181 226
rect 194 223 197 296
rect 218 286 221 306
rect 210 283 221 286
rect 210 226 213 283
rect 210 223 221 226
rect 186 193 189 206
rect 194 153 197 206
rect 218 203 221 223
rect 202 133 205 166
rect 226 163 229 463
rect 250 413 253 426
rect 250 323 253 336
rect 290 283 293 416
rect 306 406 309 416
rect 314 413 317 503
rect 322 413 325 436
rect 362 413 365 506
rect 306 403 325 406
rect 314 333 317 403
rect 362 396 365 406
rect 370 403 373 496
rect 402 493 405 526
rect 410 523 413 566
rect 418 533 421 556
rect 426 533 429 596
rect 490 593 493 616
rect 506 613 509 623
rect 434 526 437 546
rect 426 523 437 526
rect 506 523 509 606
rect 514 563 517 616
rect 522 603 525 623
rect 530 543 533 693
rect 546 676 549 806
rect 554 803 557 816
rect 562 783 565 816
rect 578 776 581 816
rect 594 783 597 816
rect 658 803 661 816
rect 666 813 669 896
rect 690 866 693 926
rect 698 896 701 933
rect 706 913 709 926
rect 810 923 813 943
rect 818 903 821 983
rect 826 923 829 966
rect 834 933 837 993
rect 858 933 861 1006
rect 698 893 709 896
rect 682 863 693 866
rect 682 813 685 863
rect 706 826 709 893
rect 706 823 717 826
rect 690 813 709 816
rect 562 773 581 776
rect 554 733 557 746
rect 562 716 565 773
rect 570 733 573 746
rect 562 713 569 716
rect 578 713 581 726
rect 594 723 597 736
rect 542 673 549 676
rect 542 616 545 673
rect 542 613 549 616
rect 538 546 541 596
rect 546 553 549 613
rect 538 543 549 546
rect 530 533 541 536
rect 426 503 429 523
rect 522 496 525 526
rect 378 396 381 416
rect 298 323 309 326
rect 322 323 325 396
rect 362 393 381 396
rect 386 353 389 406
rect 402 393 405 416
rect 418 343 421 406
rect 418 326 421 336
rect 426 333 429 496
rect 514 493 525 496
rect 514 446 517 493
rect 514 443 525 446
rect 434 333 437 426
rect 522 423 525 443
rect 530 383 533 533
rect 538 403 541 526
rect 546 406 549 536
rect 554 503 557 706
rect 566 626 569 713
rect 562 623 569 626
rect 562 583 565 623
rect 578 613 589 616
rect 570 546 573 606
rect 578 583 581 596
rect 562 543 573 546
rect 594 543 597 616
rect 602 613 605 746
rect 634 613 637 736
rect 642 733 645 796
rect 650 783 653 796
rect 666 716 669 806
rect 690 803 693 813
rect 714 806 717 823
rect 722 813 725 826
rect 818 816 821 856
rect 842 853 845 926
rect 810 813 821 816
rect 706 803 717 806
rect 682 736 685 796
rect 714 746 717 803
rect 810 793 813 813
rect 834 783 837 806
rect 858 796 861 926
rect 882 893 885 1156
rect 890 1133 893 1176
rect 898 1126 901 1193
rect 890 1123 901 1126
rect 890 886 893 1123
rect 906 1116 909 1236
rect 914 1193 917 1283
rect 930 1216 933 1293
rect 954 1266 957 1313
rect 922 1213 933 1216
rect 946 1263 957 1266
rect 914 1133 917 1146
rect 902 1113 909 1116
rect 902 1046 905 1113
rect 914 1073 917 1116
rect 922 1113 925 1213
rect 946 1196 949 1263
rect 962 1203 965 1256
rect 970 1203 973 1326
rect 978 1253 981 1336
rect 986 1323 989 1346
rect 994 1313 997 1326
rect 1026 1323 1029 1416
rect 1114 1413 1125 1416
rect 1082 1333 1085 1346
rect 1090 1333 1093 1396
rect 1114 1393 1117 1413
rect 1130 1336 1133 1526
rect 1138 1493 1141 1536
rect 1146 1523 1149 1536
rect 1154 1436 1157 1616
rect 1178 1603 1181 1626
rect 1226 1613 1237 1616
rect 1162 1443 1165 1546
rect 1170 1523 1173 1556
rect 1194 1553 1197 1606
rect 1218 1543 1221 1606
rect 1154 1433 1165 1436
rect 1138 1346 1141 1426
rect 1162 1416 1165 1433
rect 1146 1403 1149 1416
rect 1154 1413 1165 1416
rect 1170 1413 1173 1516
rect 1178 1413 1181 1526
rect 1266 1523 1269 1546
rect 1274 1513 1277 1536
rect 1282 1533 1285 1566
rect 1154 1403 1157 1413
rect 1178 1393 1181 1406
rect 1186 1403 1189 1506
rect 1138 1343 1149 1346
rect 978 1223 997 1226
rect 978 1213 981 1223
rect 986 1203 989 1216
rect 994 1213 997 1223
rect 946 1193 965 1196
rect 962 1176 965 1193
rect 898 1043 905 1046
rect 898 986 901 1043
rect 906 1013 909 1026
rect 914 1013 917 1036
rect 930 1013 933 1136
rect 938 1103 941 1176
rect 962 1173 973 1176
rect 954 1123 957 1146
rect 970 1116 973 1173
rect 962 1113 973 1116
rect 938 1013 949 1016
rect 962 1013 965 1113
rect 1002 1083 1005 1156
rect 1018 1096 1021 1196
rect 1026 1123 1029 1216
rect 1090 1203 1093 1326
rect 1098 1303 1101 1326
rect 1098 1203 1101 1296
rect 1106 1213 1109 1336
rect 1130 1333 1141 1336
rect 1130 1246 1133 1326
rect 1138 1293 1141 1333
rect 1146 1283 1149 1343
rect 1114 1243 1133 1246
rect 1114 1206 1117 1243
rect 1122 1223 1141 1226
rect 1122 1213 1133 1216
rect 1114 1203 1125 1206
rect 1042 1143 1061 1146
rect 1034 1123 1037 1136
rect 1042 1123 1045 1143
rect 1014 1093 1021 1096
rect 906 993 909 1006
rect 898 983 909 986
rect 898 906 901 926
rect 906 923 909 983
rect 922 973 925 1006
rect 938 993 941 1013
rect 946 983 949 1006
rect 898 903 905 906
rect 850 793 861 796
rect 870 883 893 886
rect 714 743 725 746
rect 682 733 693 736
rect 658 713 669 716
rect 674 613 677 716
rect 706 676 709 726
rect 714 723 717 736
rect 722 706 725 743
rect 698 673 709 676
rect 718 703 725 706
rect 730 733 741 736
rect 682 613 685 626
rect 690 613 693 636
rect 554 413 557 436
rect 562 426 565 543
rect 570 523 573 536
rect 578 533 589 536
rect 578 516 581 526
rect 570 513 581 516
rect 586 513 589 533
rect 562 423 573 426
rect 562 406 565 416
rect 546 403 565 406
rect 546 393 557 396
rect 442 326 445 346
rect 306 303 309 323
rect 234 183 237 206
rect 242 203 245 266
rect 330 263 333 326
rect 418 323 429 326
rect 250 193 253 206
rect 138 113 141 126
rect 226 123 229 156
rect 282 123 285 186
rect 330 133 333 166
rect 290 113 293 126
rect 338 123 341 216
rect 354 203 357 306
rect 370 203 373 296
rect 378 203 381 216
rect 386 186 389 206
rect 394 193 397 216
rect 402 203 405 286
rect 410 213 413 306
rect 410 186 413 206
rect 362 143 365 186
rect 386 183 413 186
rect 386 133 389 146
rect 394 123 397 156
rect 418 153 421 216
rect 426 203 429 323
rect 434 323 445 326
rect 434 303 437 323
rect 434 163 437 216
rect 442 203 445 216
rect 450 183 453 206
rect 450 133 453 146
rect 506 133 509 306
rect 530 266 533 326
rect 538 293 541 326
rect 546 323 549 336
rect 554 276 557 393
rect 562 323 565 336
rect 570 303 573 423
rect 578 416 581 506
rect 578 413 589 416
rect 578 333 581 413
rect 594 406 597 526
rect 602 413 605 556
rect 618 533 621 546
rect 610 433 613 526
rect 626 426 629 586
rect 634 523 637 606
rect 642 586 645 606
rect 642 583 653 586
rect 650 456 653 583
rect 674 523 677 546
rect 682 533 693 536
rect 642 453 653 456
rect 642 436 645 453
rect 610 423 629 426
rect 638 433 645 436
rect 610 406 613 423
rect 586 403 597 406
rect 602 403 613 406
rect 546 273 557 276
rect 530 263 541 266
rect 522 123 525 216
rect 538 213 541 263
rect 546 203 549 273
rect 554 213 557 236
rect 586 233 589 403
rect 602 386 605 403
rect 618 393 621 406
rect 594 226 597 386
rect 602 383 613 386
rect 602 343 605 383
rect 626 336 629 406
rect 638 346 641 433
rect 650 413 653 426
rect 658 413 661 436
rect 666 406 669 416
rect 650 403 669 406
rect 638 343 645 346
rect 602 313 605 336
rect 610 293 613 336
rect 622 333 629 336
rect 622 226 625 333
rect 538 133 549 136
rect 562 123 565 226
rect 586 223 605 226
rect 586 213 589 223
rect 570 123 573 206
rect 586 113 589 206
rect 594 203 597 216
rect 602 213 605 223
rect 618 223 625 226
rect 618 203 621 223
rect 634 213 637 326
rect 642 323 645 343
rect 650 266 653 403
rect 658 313 661 326
rect 642 263 653 266
rect 642 226 645 263
rect 642 223 661 226
rect 642 213 645 223
rect 650 206 653 216
rect 634 203 653 206
rect 658 186 661 223
rect 594 133 597 186
rect 654 183 661 186
rect 618 123 621 136
rect 654 126 657 183
rect 634 103 637 126
rect 642 113 645 126
rect 654 123 661 126
rect 658 103 661 123
rect 666 113 669 396
rect 674 346 677 516
rect 690 356 693 526
rect 698 523 701 673
rect 718 616 721 703
rect 706 603 709 616
rect 718 613 725 616
rect 730 613 733 733
rect 738 633 741 726
rect 762 723 765 736
rect 770 703 773 726
rect 714 583 717 596
rect 722 576 725 613
rect 714 573 725 576
rect 706 363 709 406
rect 714 403 717 573
rect 730 513 733 526
rect 738 503 741 626
rect 754 606 757 616
rect 762 613 765 626
rect 754 603 773 606
rect 794 603 797 726
rect 802 693 805 726
rect 810 713 813 736
rect 834 696 837 726
rect 826 693 837 696
rect 826 636 829 693
rect 826 633 837 636
rect 746 533 749 556
rect 754 523 757 586
rect 834 573 837 633
rect 842 566 845 696
rect 850 623 853 793
rect 870 786 873 883
rect 882 803 885 816
rect 866 783 873 786
rect 858 713 861 726
rect 866 693 869 783
rect 902 776 905 903
rect 898 773 905 776
rect 898 723 901 773
rect 914 736 917 816
rect 922 813 925 956
rect 930 916 933 966
rect 954 936 957 1006
rect 970 1003 973 1026
rect 938 933 957 936
rect 970 933 973 956
rect 938 923 941 933
rect 946 916 949 926
rect 930 913 949 916
rect 938 816 941 913
rect 962 906 965 926
rect 958 903 965 906
rect 958 846 961 903
rect 958 843 965 846
rect 962 826 965 843
rect 946 823 965 826
rect 922 773 925 806
rect 930 766 933 816
rect 938 813 957 816
rect 938 803 949 806
rect 954 796 957 813
rect 962 803 965 816
rect 954 793 965 796
rect 906 733 917 736
rect 922 763 933 766
rect 906 706 909 733
rect 898 703 909 706
rect 898 646 901 703
rect 898 643 909 646
rect 906 613 909 643
rect 914 606 917 726
rect 922 723 925 763
rect 930 713 933 736
rect 938 656 941 746
rect 962 713 965 726
rect 930 653 941 656
rect 906 603 917 606
rect 834 563 845 566
rect 778 503 781 526
rect 730 423 733 436
rect 754 403 757 426
rect 786 423 789 536
rect 794 513 797 536
rect 802 503 805 526
rect 826 516 829 526
rect 834 523 837 563
rect 842 533 845 546
rect 842 516 845 526
rect 874 523 877 596
rect 882 523 885 536
rect 826 513 845 516
rect 890 456 893 526
rect 882 453 893 456
rect 690 353 709 356
rect 674 343 685 346
rect 682 323 685 343
rect 674 296 677 316
rect 698 313 701 336
rect 674 293 685 296
rect 682 236 685 293
rect 706 276 709 353
rect 674 233 685 236
rect 698 273 709 276
rect 674 213 677 233
rect 690 203 693 216
rect 698 213 701 273
rect 706 183 709 216
rect 714 213 717 326
rect 738 306 741 366
rect 762 346 765 416
rect 882 413 885 453
rect 898 433 901 536
rect 906 523 909 603
rect 914 473 917 566
rect 898 423 917 426
rect 898 413 901 423
rect 914 416 917 423
rect 922 416 925 626
rect 930 496 933 653
rect 954 613 957 636
rect 970 633 973 926
rect 978 913 981 1036
rect 1002 1013 1005 1076
rect 1014 1026 1017 1093
rect 1014 1023 1021 1026
rect 986 923 989 966
rect 994 946 997 1006
rect 1018 963 1021 1023
rect 1026 973 1029 1116
rect 1050 1113 1053 1136
rect 1058 1133 1061 1143
rect 1082 1123 1085 1196
rect 1034 1006 1037 1016
rect 1042 1013 1045 1026
rect 1034 1003 1045 1006
rect 1018 946 1021 956
rect 994 943 1021 946
rect 994 846 997 943
rect 1002 923 1005 936
rect 1018 923 1021 936
rect 1026 916 1029 936
rect 1018 913 1029 916
rect 1034 913 1037 996
rect 1042 946 1045 1003
rect 1050 976 1053 1016
rect 1050 973 1061 976
rect 1042 943 1053 946
rect 1026 893 1029 913
rect 1042 903 1045 936
rect 1050 846 1053 943
rect 1058 923 1061 973
rect 978 843 997 846
rect 1034 843 1053 846
rect 978 813 981 843
rect 986 743 989 826
rect 978 703 981 726
rect 962 613 973 616
rect 986 613 989 736
rect 1002 676 1005 716
rect 994 673 1005 676
rect 994 613 997 673
rect 1010 636 1013 726
rect 1002 633 1013 636
rect 1002 606 1005 633
rect 946 583 949 606
rect 994 603 1005 606
rect 978 496 981 526
rect 986 523 989 536
rect 930 493 941 496
rect 730 303 741 306
rect 746 343 765 346
rect 730 236 733 303
rect 730 233 741 236
rect 722 213 733 216
rect 738 213 741 233
rect 682 133 685 156
rect 722 133 725 213
rect 674 103 677 126
rect 698 113 701 126
rect 738 123 741 206
rect 746 203 749 343
rect 754 333 765 336
rect 754 213 757 326
rect 770 313 773 326
rect 794 323 797 406
rect 810 383 813 396
rect 850 393 853 406
rect 906 386 909 416
rect 914 413 925 416
rect 922 403 925 413
rect 930 393 933 406
rect 850 356 853 386
rect 906 383 917 386
rect 850 353 869 356
rect 850 343 853 353
rect 802 323 805 336
rect 834 326 837 336
rect 858 333 861 346
rect 834 323 845 326
rect 842 236 845 323
rect 858 313 861 326
rect 842 233 853 236
rect 762 153 765 216
rect 786 143 789 216
rect 794 203 797 226
rect 802 203 805 216
rect 842 203 845 216
rect 850 213 853 233
rect 858 193 861 206
rect 866 203 869 353
rect 874 333 885 336
rect 890 333 893 376
rect 898 333 901 346
rect 874 193 877 206
rect 890 166 893 326
rect 898 313 901 326
rect 898 213 901 226
rect 882 163 893 166
rect 898 163 901 206
rect 906 183 909 356
rect 914 323 917 383
rect 938 343 941 493
rect 970 493 981 496
rect 970 436 973 493
rect 970 433 981 436
rect 978 413 981 433
rect 954 393 957 406
rect 994 353 997 603
rect 1002 343 1005 386
rect 1010 373 1013 616
rect 1018 613 1021 626
rect 1018 513 1021 526
rect 1018 393 1021 416
rect 1026 413 1029 636
rect 1034 613 1037 843
rect 1042 813 1045 836
rect 1066 813 1069 1036
rect 1090 1013 1093 1126
rect 1106 1033 1109 1146
rect 1130 1123 1133 1213
rect 1138 1026 1141 1223
rect 1146 1173 1149 1206
rect 1154 1203 1157 1306
rect 1178 1296 1181 1346
rect 1194 1333 1197 1446
rect 1250 1413 1253 1506
rect 1282 1496 1285 1526
rect 1290 1523 1293 1586
rect 1298 1513 1301 1526
rect 1322 1523 1325 1596
rect 1330 1593 1333 1606
rect 1338 1583 1341 1616
rect 1346 1573 1349 1606
rect 1354 1563 1357 1606
rect 1402 1593 1405 1616
rect 1490 1546 1493 1596
rect 1386 1526 1389 1546
rect 1482 1543 1493 1546
rect 1386 1523 1405 1526
rect 1178 1293 1189 1296
rect 1066 783 1069 806
rect 1082 803 1085 926
rect 1090 813 1093 826
rect 1090 746 1093 806
rect 1082 743 1093 746
rect 1082 726 1085 743
rect 1098 736 1101 926
rect 1106 923 1109 1026
rect 1130 1023 1141 1026
rect 1130 976 1133 1023
rect 1122 973 1133 976
rect 1114 896 1117 936
rect 1122 923 1125 973
rect 1130 933 1133 956
rect 1146 943 1149 1016
rect 1154 1013 1157 1026
rect 1114 893 1125 896
rect 1146 893 1149 926
rect 1106 813 1109 826
rect 1114 763 1117 856
rect 1122 813 1125 893
rect 1130 803 1133 826
rect 1138 813 1141 836
rect 1078 723 1085 726
rect 1090 733 1101 736
rect 1078 636 1081 723
rect 1090 646 1093 733
rect 1098 703 1101 726
rect 1122 683 1125 786
rect 1154 773 1157 1006
rect 1162 873 1165 1046
rect 1170 1013 1173 1286
rect 1186 1176 1189 1293
rect 1178 1173 1189 1176
rect 1202 1173 1205 1396
rect 1258 1383 1261 1406
rect 1210 1333 1229 1336
rect 1218 1306 1221 1326
rect 1226 1323 1229 1333
rect 1214 1303 1221 1306
rect 1214 1236 1217 1303
rect 1226 1296 1229 1316
rect 1226 1293 1237 1296
rect 1234 1246 1237 1293
rect 1226 1243 1237 1246
rect 1214 1233 1221 1236
rect 1218 1213 1221 1233
rect 1178 1053 1181 1173
rect 1202 1133 1205 1146
rect 1186 1096 1189 1126
rect 1186 1093 1197 1096
rect 1194 1036 1197 1093
rect 1186 1033 1197 1036
rect 1170 1003 1181 1006
rect 1170 953 1173 1003
rect 1178 923 1181 996
rect 1186 943 1189 1033
rect 1194 1003 1197 1016
rect 1202 943 1205 976
rect 1186 906 1189 936
rect 1194 913 1197 926
rect 1178 903 1189 906
rect 1178 826 1181 903
rect 1202 896 1205 926
rect 1194 893 1205 896
rect 1210 893 1213 1006
rect 1218 906 1221 1026
rect 1226 1003 1229 1243
rect 1234 1223 1245 1226
rect 1234 1186 1237 1223
rect 1242 1203 1245 1216
rect 1234 1183 1241 1186
rect 1238 1116 1241 1183
rect 1250 1123 1253 1216
rect 1258 1213 1261 1326
rect 1266 1213 1269 1416
rect 1274 1313 1277 1496
rect 1282 1493 1293 1496
rect 1290 1436 1293 1493
rect 1282 1433 1293 1436
rect 1282 1413 1285 1433
rect 1410 1413 1413 1536
rect 1418 1413 1421 1436
rect 1306 1333 1309 1376
rect 1314 1353 1317 1406
rect 1426 1396 1429 1536
rect 1442 1513 1445 1526
rect 1450 1493 1453 1536
rect 1482 1523 1485 1543
rect 1522 1536 1525 1606
rect 1530 1563 1533 1606
rect 1490 1513 1493 1536
rect 1522 1533 1541 1536
rect 1322 1333 1325 1396
rect 1418 1393 1429 1396
rect 1298 1213 1301 1226
rect 1266 1193 1269 1206
rect 1266 1123 1285 1126
rect 1290 1123 1293 1186
rect 1314 1183 1317 1226
rect 1238 1113 1253 1116
rect 1250 1013 1253 1113
rect 1266 1013 1269 1123
rect 1298 1046 1301 1146
rect 1290 1043 1301 1046
rect 1242 953 1245 1006
rect 1258 973 1261 1006
rect 1274 1003 1277 1016
rect 1290 1003 1293 1043
rect 1306 1036 1309 1126
rect 1314 1113 1317 1176
rect 1298 1033 1309 1036
rect 1242 933 1245 946
rect 1274 936 1277 956
rect 1234 923 1245 926
rect 1218 903 1229 906
rect 1250 903 1253 936
rect 1266 933 1277 936
rect 1178 823 1189 826
rect 1138 703 1141 726
rect 1146 713 1149 736
rect 1154 703 1157 756
rect 1162 713 1165 806
rect 1170 783 1173 796
rect 1178 733 1181 746
rect 1186 733 1189 823
rect 1194 746 1197 893
rect 1226 886 1229 903
rect 1226 883 1237 886
rect 1202 813 1205 826
rect 1210 753 1213 856
rect 1234 816 1237 883
rect 1266 846 1269 933
rect 1282 913 1285 926
rect 1266 843 1277 846
rect 1218 803 1221 816
rect 1226 813 1237 816
rect 1218 783 1221 796
rect 1226 793 1229 813
rect 1194 743 1213 746
rect 1170 693 1173 726
rect 1186 713 1189 726
rect 1194 706 1197 726
rect 1218 723 1221 776
rect 1226 733 1229 766
rect 1266 733 1269 826
rect 1274 733 1277 843
rect 1282 823 1285 896
rect 1290 816 1293 936
rect 1298 933 1301 1033
rect 1306 1003 1309 1026
rect 1314 933 1317 1046
rect 1322 983 1325 1196
rect 1330 1173 1333 1386
rect 1346 1326 1349 1356
rect 1354 1333 1357 1386
rect 1418 1383 1421 1393
rect 1434 1383 1437 1406
rect 1482 1403 1485 1416
rect 1522 1413 1525 1526
rect 1538 1416 1541 1533
rect 1554 1513 1557 1616
rect 1570 1516 1573 1606
rect 1594 1536 1597 1616
rect 1650 1563 1653 1616
rect 1578 1533 1597 1536
rect 1530 1413 1541 1416
rect 1346 1323 1357 1326
rect 1362 1323 1365 1346
rect 1338 1186 1341 1216
rect 1346 1193 1349 1206
rect 1354 1203 1357 1323
rect 1354 1186 1357 1196
rect 1338 1183 1357 1186
rect 1370 1183 1373 1336
rect 1354 1173 1357 1183
rect 1378 1133 1381 1216
rect 1386 1193 1389 1336
rect 1426 1326 1429 1346
rect 1410 1323 1429 1326
rect 1498 1323 1501 1406
rect 1514 1323 1517 1396
rect 1522 1323 1525 1406
rect 1530 1393 1533 1413
rect 1530 1333 1533 1386
rect 1562 1366 1565 1516
rect 1570 1513 1581 1516
rect 1594 1513 1597 1526
rect 1578 1436 1581 1513
rect 1570 1433 1581 1436
rect 1570 1373 1573 1433
rect 1554 1363 1565 1366
rect 1538 1333 1541 1346
rect 1410 1213 1413 1226
rect 1418 1213 1421 1236
rect 1474 1213 1477 1226
rect 1386 1133 1389 1186
rect 1330 1113 1333 1126
rect 1362 1113 1365 1126
rect 1410 1123 1413 1186
rect 1434 1173 1437 1206
rect 1330 1013 1341 1016
rect 1298 903 1301 926
rect 1282 813 1293 816
rect 1282 733 1285 813
rect 1290 726 1293 776
rect 1298 733 1301 816
rect 1314 803 1317 876
rect 1338 846 1341 1006
rect 1346 993 1349 1006
rect 1354 936 1357 1026
rect 1370 1013 1373 1036
rect 1426 1026 1429 1166
rect 1434 1143 1453 1146
rect 1434 1123 1437 1143
rect 1442 1123 1445 1136
rect 1450 1133 1453 1143
rect 1474 1123 1477 1186
rect 1490 1173 1493 1206
rect 1506 1203 1509 1306
rect 1538 1213 1541 1326
rect 1554 1176 1557 1363
rect 1578 1326 1581 1416
rect 1602 1356 1605 1406
rect 1602 1353 1613 1356
rect 1602 1333 1605 1346
rect 1570 1323 1581 1326
rect 1554 1173 1565 1176
rect 1530 1133 1533 1156
rect 1514 1113 1517 1126
rect 1554 1113 1557 1126
rect 1562 1106 1565 1173
rect 1570 1166 1573 1323
rect 1610 1316 1613 1353
rect 1626 1343 1629 1416
rect 1634 1336 1637 1526
rect 1626 1333 1637 1336
rect 1642 1333 1645 1386
rect 1690 1383 1693 1416
rect 1634 1326 1637 1333
rect 1634 1323 1645 1326
rect 1578 1296 1581 1316
rect 1602 1313 1613 1316
rect 1578 1293 1589 1296
rect 1586 1246 1589 1293
rect 1578 1243 1589 1246
rect 1578 1186 1581 1243
rect 1586 1193 1589 1216
rect 1602 1203 1605 1313
rect 1626 1196 1629 1216
rect 1578 1183 1597 1186
rect 1570 1163 1577 1166
rect 1574 1106 1577 1163
rect 1594 1156 1597 1183
rect 1602 1176 1605 1196
rect 1618 1193 1629 1196
rect 1602 1173 1613 1176
rect 1594 1153 1601 1156
rect 1554 1103 1565 1106
rect 1570 1103 1577 1106
rect 1418 1023 1429 1026
rect 1346 933 1357 936
rect 1378 933 1381 1016
rect 1418 956 1421 1023
rect 1418 953 1429 956
rect 1346 923 1349 933
rect 1338 843 1345 846
rect 1314 776 1317 796
rect 1342 776 1345 843
rect 1354 813 1357 926
rect 1426 853 1429 953
rect 1434 936 1437 1016
rect 1458 993 1461 1056
rect 1474 1013 1477 1026
rect 1434 933 1453 936
rect 1458 916 1461 936
rect 1450 913 1461 916
rect 1450 846 1453 913
rect 1450 843 1461 846
rect 1378 776 1381 836
rect 1394 813 1397 826
rect 1402 806 1405 816
rect 1314 773 1325 776
rect 1274 723 1293 726
rect 1194 703 1205 706
rect 1090 643 1097 646
rect 1034 603 1045 606
rect 1050 536 1053 636
rect 1078 633 1085 636
rect 1034 533 1053 536
rect 1034 413 1037 533
rect 1058 526 1061 536
rect 1066 533 1069 576
rect 1074 526 1077 616
rect 1082 543 1085 633
rect 1094 566 1097 643
rect 1138 603 1141 616
rect 1162 573 1165 686
rect 1178 593 1181 606
rect 1186 576 1189 696
rect 1178 573 1189 576
rect 1090 563 1097 566
rect 1042 523 1061 526
rect 1010 343 1029 346
rect 1010 333 1013 343
rect 1018 316 1021 336
rect 1010 313 1021 316
rect 914 193 917 216
rect 754 103 757 126
rect 810 123 813 136
rect 818 133 821 146
rect 882 123 885 163
rect 890 133 893 146
rect 906 133 909 146
rect 930 123 933 136
rect 938 133 941 186
rect 946 123 949 206
rect 954 123 957 236
rect 1010 213 1013 306
rect 1026 233 1029 343
rect 1034 333 1037 346
rect 1042 233 1045 516
rect 1050 406 1053 506
rect 1058 413 1061 523
rect 1066 523 1077 526
rect 1066 513 1069 523
rect 1050 403 1061 406
rect 1050 323 1053 396
rect 1066 383 1069 416
rect 1074 403 1077 436
rect 1090 423 1093 563
rect 1106 533 1109 546
rect 1098 393 1101 406
rect 1106 396 1109 416
rect 1114 403 1117 476
rect 1122 396 1125 406
rect 1106 393 1125 396
rect 1130 396 1133 416
rect 1138 413 1141 526
rect 1178 516 1181 573
rect 1202 566 1205 703
rect 1218 583 1221 706
rect 1242 623 1245 686
rect 1282 676 1285 716
rect 1298 683 1301 726
rect 1282 673 1301 676
rect 1234 603 1245 606
rect 1194 563 1205 566
rect 1194 523 1197 563
rect 1178 513 1189 516
rect 1146 416 1149 426
rect 1146 413 1173 416
rect 1130 393 1141 396
rect 1138 343 1141 393
rect 1162 346 1165 406
rect 1154 343 1165 346
rect 1146 303 1149 336
rect 1154 286 1157 343
rect 1138 283 1157 286
rect 1042 206 1045 216
rect 970 183 973 206
rect 1042 203 1053 206
rect 1042 143 1045 186
rect 1050 153 1053 203
rect 1058 113 1061 136
rect 1066 133 1069 156
rect 1074 123 1077 196
rect 1098 193 1101 206
rect 1106 203 1109 216
rect 1122 213 1125 226
rect 1114 193 1117 206
rect 1130 183 1133 216
rect 1138 203 1141 283
rect 1146 213 1149 276
rect 1154 203 1157 256
rect 1162 233 1165 326
rect 1178 313 1181 326
rect 1186 253 1189 513
rect 1218 416 1221 546
rect 1250 533 1253 616
rect 1290 606 1293 626
rect 1286 603 1293 606
rect 1210 413 1221 416
rect 1210 393 1213 413
rect 1218 363 1221 406
rect 1194 243 1197 326
rect 1202 273 1205 336
rect 1226 323 1229 416
rect 1242 413 1245 526
rect 1286 516 1289 603
rect 1298 523 1301 673
rect 1306 623 1309 756
rect 1314 733 1317 746
rect 1322 723 1325 773
rect 1338 773 1345 776
rect 1338 753 1341 773
rect 1362 733 1365 776
rect 1370 773 1381 776
rect 1394 803 1405 806
rect 1426 803 1429 816
rect 1434 813 1437 826
rect 1330 633 1333 726
rect 1354 713 1357 726
rect 1370 723 1373 773
rect 1378 713 1381 736
rect 1386 703 1389 726
rect 1394 713 1397 803
rect 1402 783 1405 796
rect 1458 786 1461 843
rect 1450 783 1461 786
rect 1402 693 1405 726
rect 1434 703 1437 726
rect 1450 696 1453 783
rect 1466 773 1469 976
rect 1474 813 1477 916
rect 1482 906 1485 996
rect 1490 923 1493 1016
rect 1514 1013 1517 1026
rect 1530 1016 1533 1046
rect 1522 1013 1533 1016
rect 1498 986 1501 1006
rect 1498 983 1509 986
rect 1506 916 1509 983
rect 1522 943 1525 1013
rect 1498 913 1509 916
rect 1482 903 1489 906
rect 1486 836 1489 903
rect 1482 833 1489 836
rect 1450 693 1461 696
rect 1362 616 1365 636
rect 1394 623 1397 656
rect 1458 623 1461 693
rect 1306 603 1309 616
rect 1358 613 1365 616
rect 1386 613 1397 616
rect 1330 553 1333 606
rect 1314 533 1317 546
rect 1346 536 1349 606
rect 1358 546 1361 613
rect 1370 573 1373 606
rect 1386 603 1397 606
rect 1358 543 1365 546
rect 1342 533 1349 536
rect 1286 513 1293 516
rect 1290 493 1293 513
rect 1242 393 1245 406
rect 1242 313 1245 336
rect 1266 323 1269 416
rect 1330 413 1333 496
rect 1342 426 1345 533
rect 1342 423 1349 426
rect 1346 406 1349 423
rect 1354 413 1357 526
rect 1362 476 1365 543
rect 1394 523 1397 596
rect 1402 583 1405 616
rect 1458 603 1461 616
rect 1482 553 1485 833
rect 1490 783 1493 816
rect 1498 776 1501 913
rect 1522 893 1525 926
rect 1506 783 1509 806
rect 1514 803 1517 826
rect 1522 813 1525 856
rect 1530 803 1533 1006
rect 1538 1003 1541 1086
rect 1554 1013 1557 1103
rect 1570 1083 1573 1103
rect 1598 1086 1601 1153
rect 1594 1083 1601 1086
rect 1546 973 1549 1006
rect 1538 923 1541 936
rect 1554 906 1557 946
rect 1546 903 1557 906
rect 1546 853 1549 903
rect 1538 813 1549 816
rect 1554 813 1557 896
rect 1498 773 1509 776
rect 1498 723 1501 736
rect 1498 586 1501 626
rect 1506 616 1509 773
rect 1562 746 1565 1006
rect 1570 1003 1573 1016
rect 1594 1013 1597 1083
rect 1522 733 1525 746
rect 1554 743 1565 746
rect 1514 653 1517 726
rect 1538 713 1541 736
rect 1554 733 1557 743
rect 1570 736 1573 956
rect 1578 833 1581 1006
rect 1602 973 1605 1006
rect 1586 933 1589 946
rect 1594 933 1597 956
rect 1610 943 1613 1173
rect 1618 1133 1621 1193
rect 1642 1133 1645 1323
rect 1690 1133 1693 1216
rect 1618 1123 1629 1126
rect 1618 1033 1621 1116
rect 1618 1003 1621 1026
rect 1586 893 1589 926
rect 1578 813 1581 826
rect 1578 793 1581 806
rect 1562 733 1573 736
rect 1578 733 1581 746
rect 1506 613 1517 616
rect 1546 613 1549 646
rect 1570 626 1573 726
rect 1586 723 1589 856
rect 1594 813 1597 926
rect 1602 906 1605 926
rect 1602 903 1609 906
rect 1606 826 1609 903
rect 1618 873 1621 926
rect 1606 823 1621 826
rect 1594 736 1597 796
rect 1602 773 1605 806
rect 1618 803 1621 823
rect 1626 813 1629 1123
rect 1634 923 1637 1036
rect 1642 913 1645 936
rect 1650 923 1653 996
rect 1658 973 1661 1016
rect 1666 1003 1669 1016
rect 1666 933 1677 936
rect 1690 923 1693 956
rect 1698 933 1701 966
rect 1634 806 1637 876
rect 1626 803 1637 806
rect 1594 733 1605 736
rect 1618 733 1621 746
rect 1594 713 1597 726
rect 1602 666 1605 733
rect 1610 706 1613 726
rect 1626 723 1629 803
rect 1666 773 1669 816
rect 1674 813 1693 816
rect 1690 793 1693 806
rect 1690 716 1693 736
rect 1682 713 1693 716
rect 1610 703 1621 706
rect 1554 623 1573 626
rect 1586 663 1605 666
rect 1490 583 1501 586
rect 1506 583 1509 606
rect 1514 593 1517 613
rect 1410 533 1413 546
rect 1362 473 1381 476
rect 1274 333 1277 366
rect 1162 203 1165 216
rect 1170 213 1173 226
rect 1178 213 1189 216
rect 1170 203 1181 206
rect 1170 143 1173 196
rect 1178 153 1181 203
rect 1274 193 1277 216
rect 1282 203 1285 226
rect 1290 213 1293 326
rect 1330 323 1333 336
rect 1338 323 1341 406
rect 1346 403 1357 406
rect 1346 333 1349 346
rect 1354 326 1357 403
rect 1378 356 1381 473
rect 1442 413 1445 526
rect 1490 523 1493 583
rect 1522 573 1525 606
rect 1538 603 1549 606
rect 1554 566 1557 586
rect 1578 573 1581 606
rect 1546 563 1557 566
rect 1506 503 1509 546
rect 1530 466 1533 526
rect 1546 486 1549 563
rect 1586 523 1589 663
rect 1618 656 1621 703
rect 1610 653 1621 656
rect 1610 623 1613 653
rect 1602 533 1605 556
rect 1626 523 1629 606
rect 1546 483 1557 486
rect 1514 463 1533 466
rect 1506 403 1509 426
rect 1514 413 1517 463
rect 1346 323 1357 326
rect 1362 353 1381 356
rect 1346 233 1349 323
rect 1362 233 1365 353
rect 1370 323 1373 336
rect 1402 333 1405 396
rect 1378 233 1381 326
rect 1394 236 1397 326
rect 1410 323 1413 396
rect 1418 243 1421 346
rect 1442 343 1445 376
rect 1394 233 1413 236
rect 1426 233 1429 326
rect 1506 323 1509 396
rect 1522 373 1525 416
rect 1538 413 1541 426
rect 1554 416 1557 483
rect 1554 413 1561 416
rect 1530 393 1533 406
rect 1546 353 1549 406
rect 1558 346 1561 413
rect 1570 396 1573 416
rect 1586 413 1589 426
rect 1602 403 1605 506
rect 1682 436 1685 713
rect 1698 626 1701 646
rect 1694 623 1701 626
rect 1694 546 1697 623
rect 1694 543 1701 546
rect 1682 433 1693 436
rect 1626 413 1629 426
rect 1690 413 1693 433
rect 1698 407 1701 543
rect 1690 404 1701 407
rect 1570 393 1581 396
rect 1082 113 1085 126
rect 1178 113 1181 136
rect 1186 133 1189 146
rect 1194 123 1197 176
rect 1202 133 1205 156
rect 1290 153 1293 206
rect 1298 173 1301 216
rect 1306 213 1309 226
rect 1210 123 1213 146
rect 1306 143 1309 206
rect 1394 193 1397 216
rect 1402 203 1405 226
rect 1410 213 1413 233
rect 1218 113 1221 126
rect 1314 113 1317 136
rect 1322 133 1325 166
rect 1330 123 1333 146
rect 1338 133 1341 156
rect 1346 123 1349 166
rect 1410 153 1413 206
rect 1418 143 1421 216
rect 1426 213 1429 226
rect 1442 143 1445 216
rect 1522 203 1525 226
rect 1530 213 1533 326
rect 1538 323 1541 336
rect 1546 333 1549 346
rect 1554 343 1561 346
rect 1514 183 1517 196
rect 1530 153 1533 206
rect 1538 203 1541 316
rect 1546 213 1549 326
rect 1554 306 1557 343
rect 1562 313 1565 326
rect 1570 323 1573 386
rect 1578 343 1581 393
rect 1690 333 1693 404
rect 1666 306 1669 326
rect 1674 313 1677 326
rect 1554 303 1573 306
rect 1666 303 1693 306
rect 1554 203 1557 246
rect 1570 206 1573 303
rect 1578 213 1581 246
rect 1586 213 1589 226
rect 1562 183 1565 206
rect 1570 203 1581 206
rect 1354 113 1357 126
rect 1450 123 1453 136
rect 1458 133 1461 146
rect 1562 143 1565 156
rect 1570 133 1573 196
rect 1578 143 1581 203
rect 1674 183 1677 196
rect 1458 113 1461 126
rect 1466 123 1477 126
rect 1586 113 1589 136
rect 1682 123 1685 246
rect 1690 203 1693 303
rect 1706 37 1726 1703
rect 1730 13 1750 1727
rect 1754 1013 1765 1016
rect 1754 813 1757 846
<< metal3 >>
rect 465 1642 510 1647
rect 329 1632 534 1637
rect 921 1632 974 1637
rect 1073 1632 1158 1637
rect 1073 1627 1078 1632
rect 505 1622 534 1627
rect 569 1622 614 1627
rect 761 1622 822 1627
rect 833 1622 1078 1627
rect 1153 1627 1158 1632
rect 1153 1622 1182 1627
rect 833 1617 838 1622
rect 457 1612 494 1617
rect 521 1612 558 1617
rect 585 1612 838 1617
rect 849 1612 910 1617
rect 1089 1612 1118 1617
rect 1201 1612 1230 1617
rect 1113 1607 1206 1612
rect 457 1602 486 1607
rect 497 1602 558 1607
rect 553 1597 558 1602
rect 641 1602 710 1607
rect 641 1597 646 1602
rect 289 1592 334 1597
rect 449 1592 534 1597
rect 553 1592 646 1597
rect 665 1592 774 1597
rect 801 1592 846 1597
rect 897 1592 950 1597
rect 977 1592 1102 1597
rect 1329 1592 1406 1597
rect 321 1582 358 1587
rect 473 1582 534 1587
rect 1121 1582 1214 1587
rect 1289 1582 1342 1587
rect 1121 1577 1126 1582
rect 201 1572 286 1577
rect 961 1572 1126 1577
rect 1209 1577 1214 1582
rect 1209 1572 1350 1577
rect 377 1562 430 1567
rect 1281 1562 1654 1567
rect 417 1547 422 1557
rect 945 1552 974 1557
rect 969 1547 974 1552
rect 1057 1552 1198 1557
rect 1057 1547 1062 1552
rect 361 1542 446 1547
rect 625 1542 670 1547
rect 697 1542 734 1547
rect 769 1542 902 1547
rect 969 1542 1062 1547
rect 1161 1542 1222 1547
rect 0 1532 86 1537
rect 105 1527 110 1537
rect 473 1532 670 1537
rect 785 1532 878 1537
rect 1081 1532 1150 1537
rect 105 1522 126 1527
rect 281 1522 334 1527
rect 457 1522 494 1527
rect 649 1522 750 1527
rect 809 1522 878 1527
rect 1249 1522 1270 1527
rect 1281 1522 1326 1527
rect 129 1512 190 1517
rect 305 1512 342 1517
rect 521 1512 566 1517
rect 649 1512 678 1517
rect 721 1512 766 1517
rect 833 1512 894 1517
rect 1105 1512 1174 1517
rect 81 1502 158 1507
rect 177 1502 278 1507
rect 321 1502 358 1507
rect 449 1502 550 1507
rect 761 1502 790 1507
rect 785 1497 790 1502
rect 881 1502 910 1507
rect 1121 1502 1190 1507
rect 1249 1502 1254 1522
rect 1273 1512 1302 1517
rect 1441 1512 1494 1517
rect 1553 1512 1598 1517
rect 881 1497 886 1502
rect 425 1492 534 1497
rect 785 1492 886 1497
rect 1137 1492 1166 1497
rect 1161 1487 1166 1492
rect 1249 1492 1454 1497
rect 1249 1487 1254 1492
rect 1161 1482 1254 1487
rect 217 1462 350 1467
rect 217 1457 222 1462
rect 193 1452 222 1457
rect 345 1457 350 1462
rect 345 1452 566 1457
rect 129 1442 158 1447
rect 601 1442 790 1447
rect 849 1442 1142 1447
rect 1161 1442 1198 1447
rect 177 1437 246 1442
rect 1137 1437 1142 1442
rect 105 1432 182 1437
rect 241 1432 334 1437
rect 793 1432 918 1437
rect 929 1432 1006 1437
rect 1137 1432 1422 1437
rect 913 1427 918 1432
rect 161 1422 230 1427
rect 225 1417 230 1422
rect 313 1422 342 1427
rect 377 1422 454 1427
rect 745 1422 782 1427
rect 913 1422 942 1427
rect 313 1417 318 1422
rect 169 1412 206 1417
rect 225 1412 318 1417
rect 609 1412 758 1417
rect 857 1412 910 1417
rect 1145 1412 1182 1417
rect 489 1402 518 1407
rect 1481 1402 1526 1407
rect 137 1392 166 1397
rect 993 1392 1094 1397
rect 1177 1392 1206 1397
rect 1513 1392 1534 1397
rect 321 1382 382 1387
rect 425 1382 686 1387
rect 1257 1382 1422 1387
rect 1433 1382 1694 1387
rect 1305 1372 1374 1377
rect 1369 1367 1374 1372
rect 1545 1372 1606 1377
rect 1545 1367 1550 1372
rect 593 1362 678 1367
rect 1369 1362 1550 1367
rect 249 1352 310 1357
rect 1313 1352 1350 1357
rect 145 1342 182 1347
rect 273 1342 358 1347
rect 617 1342 758 1347
rect 777 1342 878 1347
rect 953 1342 990 1347
rect 1177 1342 1310 1347
rect 1361 1342 1542 1347
rect 1601 1342 1630 1347
rect 89 1332 254 1337
rect 497 1332 518 1337
rect 945 1332 966 1337
rect 1081 1332 1110 1337
rect 241 1322 342 1327
rect 1025 1322 1094 1327
rect 1497 1317 1502 1327
rect 113 1312 190 1317
rect 289 1312 326 1317
rect 521 1312 694 1317
rect 961 1312 998 1317
rect 1225 1312 1278 1317
rect 1497 1312 1510 1317
rect 97 1302 134 1307
rect 233 1302 302 1307
rect 393 1302 430 1307
rect 513 1302 558 1307
rect 977 1302 1006 1307
rect 1001 1297 1006 1302
rect 1073 1302 1158 1307
rect 1505 1302 1510 1312
rect 1073 1297 1078 1302
rect 289 1292 310 1297
rect 1001 1292 1078 1297
rect 1097 1292 1142 1297
rect 265 1282 406 1287
rect 1145 1282 1174 1287
rect 785 1262 926 1267
rect 785 1257 790 1262
rect 625 1252 790 1257
rect 625 1247 630 1252
rect 281 1237 286 1247
rect 313 1242 366 1247
rect 377 1242 446 1247
rect 601 1242 630 1247
rect 921 1247 926 1262
rect 961 1252 982 1257
rect 1281 1252 1486 1257
rect 1281 1247 1286 1252
rect 921 1242 1286 1247
rect 1481 1247 1486 1252
rect 1481 1242 1510 1247
rect 249 1232 318 1237
rect 801 1232 910 1237
rect 1353 1232 1422 1237
rect 225 1222 262 1227
rect 281 1222 350 1227
rect 497 1222 542 1227
rect 569 1222 678 1227
rect 713 1222 758 1227
rect 673 1217 678 1222
rect 337 1212 374 1217
rect 529 1212 566 1217
rect 673 1212 742 1217
rect 0 1202 86 1207
rect 185 1202 318 1207
rect 657 1202 694 1207
rect 185 1197 190 1202
rect 105 1192 190 1197
rect 313 1197 318 1202
rect 313 1192 758 1197
rect 201 1182 350 1187
rect 801 1182 806 1227
rect 1297 1222 1318 1227
rect 849 1182 854 1217
rect 1025 1212 1110 1217
rect 1241 1212 1262 1217
rect 969 1202 990 1207
rect 913 1192 1022 1197
rect 1265 1192 1326 1197
rect 1345 1192 1390 1197
rect 1041 1182 1126 1187
rect 1289 1182 1318 1187
rect 1369 1182 1390 1187
rect 1409 1182 1414 1227
rect 1473 1182 1478 1227
rect 1585 1192 1606 1197
rect 561 1177 630 1182
rect 1041 1177 1046 1182
rect 249 1172 350 1177
rect 457 1172 566 1177
rect 625 1172 750 1177
rect 825 1172 878 1177
rect 889 1172 1046 1177
rect 1121 1177 1126 1182
rect 1513 1177 1670 1182
rect 1121 1172 1302 1177
rect 1313 1172 1334 1177
rect 1353 1172 1518 1177
rect 1665 1172 1694 1177
rect 1297 1167 1302 1172
rect 193 1162 238 1167
rect 329 1162 358 1167
rect 457 1162 486 1167
rect 481 1157 486 1162
rect 577 1162 606 1167
rect 769 1162 886 1167
rect 1297 1162 1558 1167
rect 577 1157 582 1162
rect 1089 1157 1158 1162
rect 1553 1157 1558 1162
rect 1617 1162 1646 1167
rect 1617 1157 1622 1162
rect 305 1152 334 1157
rect 481 1152 582 1157
rect 817 1152 886 1157
rect 1001 1152 1094 1157
rect 1153 1152 1182 1157
rect 1217 1152 1414 1157
rect 1217 1147 1222 1152
rect 1409 1147 1414 1152
rect 1505 1152 1534 1157
rect 1553 1152 1622 1157
rect 1505 1147 1510 1152
rect 105 1142 142 1147
rect 281 1142 326 1147
rect 737 1142 822 1147
rect 913 1142 958 1147
rect 1105 1142 1222 1147
rect 1297 1142 1390 1147
rect 1409 1142 1510 1147
rect 369 1132 414 1137
rect 537 1132 614 1137
rect 753 1132 934 1137
rect 305 1122 462 1127
rect 809 1122 1038 1127
rect 1313 1122 1446 1127
rect 89 1112 134 1117
rect 217 1112 342 1117
rect 873 1112 926 1117
rect 1025 1112 1318 1117
rect 1329 1112 1366 1117
rect 1513 1112 1558 1117
rect 737 1102 942 1107
rect 361 1092 582 1097
rect 361 1087 366 1092
rect 137 1082 366 1087
rect 577 1087 582 1092
rect 577 1082 734 1087
rect 729 1077 734 1082
rect 889 1082 1006 1087
rect 1537 1082 1574 1087
rect 889 1077 894 1082
rect 729 1072 894 1077
rect 913 1072 1006 1077
rect 1297 1072 1438 1077
rect 225 1062 566 1067
rect 1297 1057 1302 1072
rect 137 1052 206 1057
rect 529 1052 582 1057
rect 841 1052 998 1057
rect 137 1047 142 1052
rect 201 1047 510 1052
rect 841 1047 846 1052
rect 113 1042 142 1047
rect 505 1042 574 1047
rect 817 1042 846 1047
rect 993 1047 998 1052
rect 1025 1052 1142 1057
rect 1177 1052 1302 1057
rect 1433 1057 1438 1072
rect 1433 1052 1462 1057
rect 1553 1052 1767 1057
rect 1025 1047 1030 1052
rect 993 1042 1030 1047
rect 1137 1047 1142 1052
rect 1553 1047 1558 1052
rect 1137 1042 1166 1047
rect 1313 1042 1558 1047
rect 0 1032 70 1037
rect 161 1032 582 1037
rect 793 1032 918 1037
rect 929 1032 982 1037
rect 1065 1032 1110 1037
rect 1369 1032 1767 1037
rect 65 1027 70 1032
rect 65 1022 182 1027
rect 201 1022 246 1027
rect 321 1022 358 1027
rect 409 1022 454 1027
rect 601 1022 694 1027
rect 905 1022 974 1027
rect 1041 1022 1222 1027
rect 1265 1022 1310 1027
rect 1353 1022 1478 1027
rect 1513 1022 1622 1027
rect 0 1012 30 1017
rect 137 1012 166 1017
rect 25 1007 142 1012
rect 177 1007 182 1022
rect 601 1017 606 1022
rect 257 1012 366 1017
rect 473 1012 502 1017
rect 545 1012 606 1017
rect 689 1017 694 1022
rect 689 1012 742 1017
rect 865 1012 894 1017
rect 1009 1012 1038 1017
rect 1337 1012 1366 1017
rect 1505 1012 1670 1017
rect 1753 1012 1767 1017
rect 257 1007 262 1012
rect 889 1007 1014 1012
rect 1361 1007 1510 1012
rect 177 1002 262 1007
rect 481 1002 678 1007
rect 745 1002 862 1007
rect 1049 1002 1278 1007
rect 1529 1002 1574 1007
rect 0 992 94 997
rect 281 992 510 997
rect 905 992 1038 997
rect 1177 992 1350 997
rect 1457 992 1486 997
rect 1649 992 1767 997
rect 537 987 814 992
rect 81 982 350 987
rect 513 982 542 987
rect 809 982 926 987
rect 945 982 1382 987
rect 369 977 494 982
rect 273 972 374 977
rect 489 972 902 977
rect 921 972 1030 977
rect 1201 972 1286 977
rect 1393 972 1606 977
rect 1657 972 1767 977
rect 897 967 902 972
rect 1281 967 1398 972
rect 345 962 678 967
rect 769 962 830 967
rect 897 962 934 967
rect 985 962 1022 967
rect 1553 962 1702 967
rect 233 952 334 957
rect 449 952 550 957
rect 329 947 454 952
rect 673 947 678 962
rect 1553 957 1558 962
rect 689 952 798 957
rect 817 952 974 957
rect 1017 952 1206 957
rect 1241 952 1342 957
rect 817 947 822 952
rect 1337 947 1342 952
rect 1497 952 1558 957
rect 1569 952 1598 957
rect 1689 952 1767 957
rect 1497 947 1502 952
rect 473 942 534 947
rect 673 942 822 947
rect 857 942 1070 947
rect 1185 942 1246 947
rect 1337 942 1502 947
rect 1521 942 1558 947
rect 1585 942 1614 947
rect 129 932 278 937
rect 329 932 1006 937
rect 1249 932 1318 937
rect 1537 932 1670 937
rect 1697 932 1767 937
rect 129 927 134 932
rect 0 922 70 927
rect 97 922 134 927
rect 337 922 366 927
rect 457 922 518 927
rect 617 922 734 927
rect 833 922 862 927
rect 905 922 974 927
rect 1017 922 1238 927
rect 1593 922 1638 927
rect 65 912 70 922
rect 361 917 462 922
rect 729 917 838 922
rect 481 912 590 917
rect 681 912 710 917
rect 977 912 1022 917
rect 1033 912 1270 917
rect 1281 912 1646 917
rect 1665 912 1767 917
rect 1265 907 1270 912
rect 1665 907 1670 912
rect 0 902 30 907
rect 25 897 30 902
rect 129 902 158 907
rect 345 902 478 907
rect 489 902 518 907
rect 129 897 134 902
rect 25 892 134 897
rect 513 897 518 902
rect 641 902 910 907
rect 641 897 646 902
rect 905 897 910 902
rect 1001 902 1046 907
rect 1145 902 1254 907
rect 1265 902 1302 907
rect 1561 902 1670 907
rect 1001 897 1006 902
rect 513 892 646 897
rect 665 892 694 897
rect 689 887 694 892
rect 857 892 886 897
rect 905 892 1006 897
rect 1025 892 1150 897
rect 1209 892 1286 897
rect 1521 892 1590 897
rect 1681 892 1767 897
rect 857 887 862 892
rect 1601 887 1686 892
rect 689 882 862 887
rect 1153 882 1606 887
rect 1161 872 1190 877
rect 1289 872 1318 877
rect 1545 872 1622 877
rect 1633 872 1767 877
rect 1185 867 1294 872
rect 377 862 494 867
rect 1025 862 1094 867
rect 1025 857 1030 862
rect 193 852 230 857
rect 817 852 846 857
rect 921 852 1030 857
rect 1089 857 1094 862
rect 1337 862 1406 867
rect 1337 857 1342 862
rect 1089 852 1118 857
rect 1209 852 1342 857
rect 1401 857 1406 862
rect 1609 857 1742 862
rect 1401 852 1430 857
rect 1521 852 1550 857
rect 1585 852 1614 857
rect 1737 852 1767 857
rect 209 842 278 847
rect 521 842 598 847
rect 1121 842 1198 847
rect 1353 842 1758 847
rect 89 832 214 837
rect 65 817 70 827
rect 345 822 390 827
rect 0 812 70 817
rect 361 812 390 817
rect 169 802 342 807
rect 385 802 390 812
rect 401 797 406 817
rect 537 812 582 817
rect 593 812 598 842
rect 1193 837 1358 842
rect 1041 832 1142 837
rect 1377 832 1606 837
rect 1737 832 1767 837
rect 1601 827 1742 832
rect 721 817 726 827
rect 985 822 1094 827
rect 1105 822 1134 827
rect 1201 822 1270 827
rect 1393 822 1518 827
rect 1529 822 1582 827
rect 657 812 726 817
rect 921 812 966 817
rect 1065 812 1094 817
rect 1545 812 1694 817
rect 1753 812 1767 817
rect 537 802 646 807
rect 881 802 942 807
rect 1089 802 1094 812
rect 1161 802 1222 807
rect 1265 802 1430 807
rect 1489 802 1534 807
rect 0 792 110 797
rect 353 792 406 797
rect 417 792 542 797
rect 641 792 646 802
rect 961 792 1318 797
rect 1577 792 1598 797
rect 1689 792 1767 797
rect 417 787 422 792
rect 361 782 422 787
rect 521 782 566 787
rect 593 782 654 787
rect 833 782 1126 787
rect 1169 782 1494 787
rect 1505 782 1630 787
rect 177 772 254 777
rect 273 772 382 777
rect 401 772 430 777
rect 921 772 950 777
rect 1153 772 1222 777
rect 1289 772 1366 777
rect 1465 772 1494 777
rect 945 767 950 772
rect 1489 767 1494 772
rect 1577 772 1606 777
rect 1665 772 1767 777
rect 1577 767 1582 772
rect 217 762 238 767
rect 329 762 382 767
rect 441 762 550 767
rect 945 762 1078 767
rect 1113 762 1230 767
rect 1489 762 1582 767
rect 377 757 446 762
rect 1073 757 1078 762
rect 225 752 270 757
rect 153 742 198 747
rect 353 727 358 757
rect 1073 752 1214 757
rect 1225 752 1294 757
rect 1305 752 1342 757
rect 409 742 502 747
rect 521 742 574 747
rect 937 742 990 747
rect 1177 742 1318 747
rect 1361 742 1622 747
rect 401 732 526 737
rect 553 732 598 737
rect 689 732 718 737
rect 1169 732 1190 737
rect 1169 727 1174 732
rect 353 722 398 727
rect 497 722 542 727
rect 633 722 766 727
rect 1169 722 1198 727
rect 289 712 406 717
rect 577 712 662 717
rect 673 712 814 717
rect 857 712 934 717
rect 961 712 1014 717
rect 1145 712 1190 717
rect 1281 712 1286 737
rect 257 702 310 707
rect 305 697 310 702
rect 417 702 558 707
rect 769 702 894 707
rect 417 697 422 702
rect 889 697 894 702
rect 953 702 982 707
rect 1097 702 1142 707
rect 1153 702 1222 707
rect 953 697 958 702
rect 1297 697 1302 737
rect 1321 732 1406 737
rect 1401 727 1406 732
rect 1473 732 1542 737
rect 1569 732 1694 737
rect 1473 727 1478 732
rect 1401 722 1478 727
rect 1353 712 1382 717
rect 1537 712 1598 717
rect 1385 702 1438 707
rect 305 692 422 697
rect 737 692 870 697
rect 889 692 958 697
rect 1009 692 1174 697
rect 1185 692 1302 697
rect 1329 692 1406 697
rect 1121 682 1166 687
rect 1241 682 1302 687
rect 0 672 110 677
rect 393 662 518 667
rect 1417 662 1494 667
rect 1417 657 1422 662
rect 1009 652 1374 657
rect 1393 652 1422 657
rect 1489 657 1494 662
rect 1489 652 1518 657
rect 1009 647 1014 652
rect 985 642 1014 647
rect 1369 647 1374 652
rect 1369 642 1702 647
rect 1217 637 1310 642
rect 121 632 198 637
rect 689 632 742 637
rect 953 632 1030 637
rect 1049 632 1222 637
rect 1305 632 1366 637
rect 65 617 70 627
rect 217 622 326 627
rect 681 622 854 627
rect 905 622 926 627
rect 993 622 1062 627
rect 1289 622 1310 627
rect 1457 622 1502 627
rect 993 617 998 622
rect 1057 617 1238 622
rect 0 612 70 617
rect 105 612 134 617
rect 185 612 366 617
rect 585 612 710 617
rect 969 612 998 617
rect 1009 612 1038 617
rect 1233 612 1390 617
rect 201 602 262 607
rect 273 602 294 607
rect 313 602 342 607
rect 793 602 1038 607
rect 1137 602 1238 607
rect 1305 602 1390 607
rect 1457 602 1542 607
rect 289 597 294 602
rect 89 592 134 597
rect 289 592 366 597
rect 425 592 494 597
rect 1073 592 1182 597
rect 1249 592 1350 597
rect 1393 592 1518 597
rect 817 587 926 592
rect 537 582 630 587
rect 713 582 822 587
rect 921 582 950 587
rect 1217 582 1374 587
rect 1401 582 1558 587
rect 401 577 510 582
rect 377 572 406 577
rect 505 572 534 577
rect 833 572 1070 577
rect 1161 572 1206 577
rect 529 567 766 572
rect 1201 567 1206 572
rect 1305 572 1334 577
rect 1369 572 1582 577
rect 1305 567 1310 572
rect 409 562 518 567
rect 761 562 822 567
rect 889 562 918 567
rect 1201 562 1310 567
rect 817 557 894 562
rect 1353 557 1462 562
rect 353 552 510 557
rect 545 552 606 557
rect 633 552 750 557
rect 1329 552 1358 557
rect 1457 552 1606 557
rect 529 537 534 547
rect 593 542 622 547
rect 673 542 846 547
rect 1081 542 1510 547
rect 529 532 550 537
rect 569 532 686 537
rect 785 532 886 537
rect 1057 532 1094 537
rect 0 522 70 527
rect 65 512 70 522
rect 129 502 134 527
rect 337 522 382 527
rect 505 522 598 527
rect 881 522 990 527
rect 337 497 342 522
rect 881 517 886 522
rect 1089 517 1094 532
rect 1225 532 1254 537
rect 1225 517 1230 532
rect 545 512 574 517
rect 585 512 678 517
rect 729 512 798 517
rect 841 512 886 517
rect 1017 512 1070 517
rect 1089 512 1230 517
rect 361 502 430 507
rect 553 502 582 507
rect 689 502 742 507
rect 777 502 830 507
rect 825 497 830 502
rect 889 502 1054 507
rect 1505 502 1606 507
rect 889 497 894 502
rect 337 492 374 497
rect 401 492 430 497
rect 825 492 894 497
rect 1289 492 1334 497
rect 0 472 158 477
rect 193 472 230 477
rect 913 472 1118 477
rect 185 442 302 447
rect 185 437 190 442
rect 137 432 190 437
rect 297 437 302 442
rect 921 442 1054 447
rect 921 437 926 442
rect 297 432 326 437
rect 553 432 806 437
rect 897 432 926 437
rect 1049 437 1054 442
rect 1049 432 1078 437
rect 801 427 806 432
rect 201 422 254 427
rect 433 422 526 427
rect 649 422 718 427
rect 753 422 790 427
rect 801 422 1030 427
rect 1089 422 1150 427
rect 1505 422 1542 427
rect 1585 422 1630 427
rect 289 412 374 417
rect 1113 412 1190 417
rect 1225 412 1246 417
rect 665 402 758 407
rect 921 402 958 407
rect 321 392 406 397
rect 617 392 670 397
rect 849 392 934 397
rect 1017 392 1054 397
rect 1097 392 1166 397
rect 1209 392 1246 397
rect 1401 392 1534 397
rect 313 382 342 387
rect 337 377 342 382
rect 417 382 598 387
rect 609 382 854 387
rect 1001 382 1070 387
rect 417 377 422 382
rect 337 372 422 377
rect 889 372 1014 377
rect 1441 372 1526 377
rect 705 362 742 367
rect 777 362 1278 367
rect 777 357 782 362
rect 97 352 142 357
rect 385 352 694 357
rect 753 352 782 357
rect 905 352 998 357
rect 1521 352 1550 357
rect 129 342 158 347
rect 177 332 254 337
rect 417 332 422 352
rect 689 347 758 352
rect 1521 347 1526 352
rect 793 342 862 347
rect 897 342 1038 347
rect 1185 342 1526 347
rect 1545 342 1694 347
rect 561 332 582 337
rect 761 332 806 337
rect 873 332 902 337
rect 1049 332 1174 337
rect 1305 332 1398 337
rect 897 327 1054 332
rect 1169 327 1310 332
rect 1393 327 1398 332
rect 1481 332 1542 337
rect 1481 327 1486 332
rect 0 322 134 327
rect 129 312 134 322
rect 0 302 86 307
rect 161 302 166 327
rect 209 322 638 327
rect 1329 322 1374 327
rect 1393 322 1486 327
rect 1505 317 1510 327
rect 1545 322 1574 327
rect 601 312 678 317
rect 697 312 774 317
rect 857 312 1014 317
rect 1177 312 1246 317
rect 1505 312 1542 317
rect 1561 312 1678 317
rect 193 302 222 307
rect 305 302 358 307
rect 409 302 438 307
rect 505 302 574 307
rect 1009 302 1150 307
rect 105 292 198 297
rect 369 292 614 297
rect 289 282 406 287
rect 0 272 182 277
rect 1145 272 1206 277
rect 241 262 334 267
rect 1153 252 1190 257
rect 1441 252 1534 257
rect 1441 247 1446 252
rect 1193 242 1222 247
rect 1417 242 1446 247
rect 1529 247 1534 252
rect 1529 242 1558 247
rect 1577 242 1686 247
rect 553 232 590 237
rect 953 232 1030 237
rect 0 222 126 227
rect 137 222 182 227
rect 561 222 638 227
rect 697 222 758 227
rect 793 222 902 227
rect 273 212 358 217
rect 401 212 446 217
rect 689 212 718 217
rect 737 212 806 217
rect 865 212 918 217
rect 1041 212 1046 237
rect 1161 232 1206 237
rect 1121 222 1174 227
rect 1105 212 1182 217
rect 273 207 278 212
rect 249 202 278 207
rect 353 207 358 212
rect 353 202 382 207
rect 545 202 598 207
rect 617 202 742 207
rect 841 202 878 207
rect 1097 202 1166 207
rect 897 197 990 202
rect 1201 197 1206 232
rect 1217 217 1222 242
rect 1281 222 1310 227
rect 1217 212 1278 217
rect 1289 207 1294 217
rect 1289 202 1310 207
rect 1345 197 1350 237
rect 185 192 398 197
rect 857 192 902 197
rect 985 192 1118 197
rect 1169 192 1206 197
rect 1289 192 1350 197
rect 233 182 526 187
rect 593 182 710 187
rect 905 182 974 187
rect 1041 182 1134 187
rect 1193 172 1302 177
rect 1033 167 1174 172
rect 201 162 230 167
rect 329 162 438 167
rect 897 162 1038 167
rect 1169 162 1350 167
rect 1361 157 1366 237
rect 1377 217 1382 237
rect 1425 232 1462 237
rect 1401 222 1430 227
rect 1377 212 1398 217
rect 1409 212 1446 217
rect 1457 187 1462 232
rect 1521 222 1590 227
rect 1529 212 1574 217
rect 1569 192 1574 212
rect 1457 182 1518 187
rect 1561 182 1678 187
rect 193 152 230 157
rect 393 152 422 157
rect 681 152 766 157
rect 1049 152 1182 157
rect 1201 152 1294 157
rect 1337 152 1414 157
rect 1529 152 1566 157
rect 385 142 454 147
rect 721 142 822 147
rect 889 142 1038 147
rect 1137 142 1214 147
rect 1329 142 1422 147
rect 1457 142 1582 147
rect 1033 137 1142 142
rect 545 132 622 137
rect 809 132 910 137
rect 1161 127 1238 132
rect 929 122 958 127
rect 953 117 958 122
rect 1033 122 1166 127
rect 1233 122 1382 127
rect 1449 122 1470 127
rect 1033 117 1038 122
rect 1377 117 1382 122
rect 137 112 294 117
rect 585 112 646 117
rect 665 112 702 117
rect 953 112 1038 117
rect 1057 112 1086 117
rect 1177 112 1222 117
rect 1313 112 1358 117
rect 1377 112 1590 117
rect 633 102 758 107
use CORDIC_TOP_VIA1  CORDIC_TOP_VIA1_0
timestamp 1683038052
transform 1 0 24 0 1 1717
box -10 -10 10 10
use CORDIC_TOP_VIA1  CORDIC_TOP_VIA1_1
timestamp 1683038052
transform 1 0 1740 0 1 1717
box -10 -10 10 10
use CORDIC_TOP_VIA1  CORDIC_TOP_VIA1_2
timestamp 1683038052
transform 1 0 48 0 1 1693
box -10 -10 10 10
use CORDIC_TOP_VIA1  CORDIC_TOP_VIA1_3
timestamp 1683038052
transform 1 0 1716 0 1 1693
box -10 -10 10 10
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_0
timestamp 1683038052
transform 1 0 24 0 1 1670
box -10 -3 10 3
use M2_M1  M2_M1_14
timestamp 1683038052
transform 1 0 148 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_43
timestamp 1683038052
transform 1 0 108 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1683038052
transform 1 0 204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1683038052
transform 1 0 212 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1683038052
transform 1 0 268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1683038052
transform 1 0 292 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_29
timestamp 1683038052
transform 1 0 292 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1683038052
transform 1 0 316 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1683038052
transform 1 0 332 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_18
timestamp 1683038052
transform 1 0 356 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1683038052
transform 1 0 332 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_31
timestamp 1683038052
transform 1 0 332 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1683038052
transform 1 0 324 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_46
timestamp 1683038052
transform 1 0 356 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_3
timestamp 1683038052
transform 1 0 420 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_0
timestamp 1683038052
transform 1 0 468 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_0
timestamp 1683038052
transform 1 0 452 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_4
timestamp 1683038052
transform 1 0 460 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1683038052
transform 1 0 444 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_14
timestamp 1683038052
transform 1 0 460 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1683038052
transform 1 0 508 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_1
timestamp 1683038052
transform 1 0 508 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_3
timestamp 1683038052
transform 1 0 532 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_5
timestamp 1683038052
transform 1 0 492 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1683038052
transform 1 0 500 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_6
timestamp 1683038052
transform 1 0 508 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_7
timestamp 1683038052
transform 1 0 524 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_7
timestamp 1683038052
transform 1 0 532 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_20
timestamp 1683038052
transform 1 0 476 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_15
timestamp 1683038052
transform 1 0 492 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_21
timestamp 1683038052
transform 1 0 508 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_16
timestamp 1683038052
transform 1 0 524 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_8
timestamp 1683038052
transform 1 0 556 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1683038052
transform 1 0 532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_23
timestamp 1683038052
transform 1 0 540 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_25
timestamp 1683038052
transform 1 0 460 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_46
timestamp 1683038052
transform 1 0 468 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_26
timestamp 1683038052
transform 1 0 484 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_47
timestamp 1683038052
transform 1 0 492 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_27
timestamp 1683038052
transform 1 0 500 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_48
timestamp 1683038052
transform 1 0 532 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_32
timestamp 1683038052
transform 1 0 452 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1683038052
transform 1 0 476 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1683038052
transform 1 0 532 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_48
timestamp 1683038052
transform 1 0 532 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1683038052
transform 1 0 556 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1683038052
transform 1 0 572 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_49
timestamp 1683038052
transform 1 0 572 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_9
timestamp 1683038052
transform 1 0 612 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1683038052
transform 1 0 588 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1683038052
transform 1 0 764 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_24
timestamp 1683038052
transform 1 0 612 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1683038052
transform 1 0 668 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1683038052
transform 1 0 588 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_19
timestamp 1683038052
transform 1 0 684 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_26
timestamp 1683038052
transform 1 0 708 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1683038052
transform 1 0 764 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1683038052
transform 1 0 684 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_28
timestamp 1683038052
transform 1 0 708 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1683038052
transform 1 0 668 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_52
timestamp 1683038052
transform 1 0 772 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_35
timestamp 1683038052
transform 1 0 772 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_2
timestamp 1683038052
transform 1 0 820 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_9
timestamp 1683038052
transform 1 0 812 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_11
timestamp 1683038052
transform 1 0 820 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_28
timestamp 1683038052
transform 1 0 804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1683038052
transform 1 0 820 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_36
timestamp 1683038052
transform 1 0 804 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_10
timestamp 1683038052
transform 1 0 852 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_12
timestamp 1683038052
transform 1 0 860 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1683038052
transform 1 0 852 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_53
timestamp 1683038052
transform 1 0 844 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_37
timestamp 1683038052
transform 1 0 844 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_11
timestamp 1683038052
transform 1 0 884 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1683038052
transform 1 0 868 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_21
timestamp 1683038052
transform 1 0 884 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_31
timestamp 1683038052
transform 1 0 900 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_22
timestamp 1683038052
transform 1 0 908 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4
timestamp 1683038052
transform 1 0 924 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_32
timestamp 1683038052
transform 1 0 916 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1683038052
transform 1 0 908 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_38
timestamp 1683038052
transform 1 0 900 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_12
timestamp 1683038052
transform 1 0 932 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_5
timestamp 1683038052
transform 1 0 972 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_13
timestamp 1683038052
transform 1 0 964 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1683038052
transform 1 0 964 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_39
timestamp 1683038052
transform 1 0 948 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1683038052
transform 1 0 1180 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_33
timestamp 1683038052
transform 1 0 988 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1683038052
transform 1 0 996 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1683038052
transform 1 0 980 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_23
timestamp 1683038052
transform 1 0 1092 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_35
timestamp 1683038052
transform 1 0 1100 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1683038052
transform 1 0 1156 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1683038052
transform 1 0 1092 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1683038052
transform 1 0 1180 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_40
timestamp 1683038052
transform 1 0 980 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1683038052
transform 1 0 1020 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_67
timestamp 1683038052
transform 1 0 1084 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_42
timestamp 1683038052
transform 1 0 1100 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_59
timestamp 1683038052
transform 1 0 1196 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_24
timestamp 1683038052
transform 1 0 1228 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_37
timestamp 1683038052
transform 1 0 1236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1683038052
transform 1 0 1340 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_60
timestamp 1683038052
transform 1 0 1220 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1683038052
transform 1 0 1332 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1683038052
transform 1 0 1324 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_43
timestamp 1683038052
transform 1 0 1332 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_62
timestamp 1683038052
transform 1 0 1348 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1683038052
transform 1 0 1356 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_49
timestamp 1683038052
transform 1 0 1292 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_50
timestamp 1683038052
transform 1 0 1340 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_39
timestamp 1683038052
transform 1 0 1404 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_44
timestamp 1683038052
transform 1 0 1404 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_69
timestamp 1683038052
transform 1 0 1492 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1683038052
transform 1 0 1524 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_65
timestamp 1683038052
transform 1 0 1532 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1683038052
transform 1 0 1556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1683038052
transform 1 0 1596 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1683038052
transform 1 0 1652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1683038052
transform 1 0 1572 0 1 1605
box -2 -2 2 2
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_1
timestamp 1683038052
transform 1 0 1740 0 1 1670
box -10 -3 10 3
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_2
timestamp 1683038052
transform 1 0 48 0 1 1570
box -10 -3 10 3
use FILL  FILL_0
timestamp 1683038052
transform 1 0 72 0 1 1570
box -8 -3 16 105
use FILL  FILL_1
timestamp 1683038052
transform 1 0 80 0 1 1570
box -8 -3 16 105
use FILL  FILL_2
timestamp 1683038052
transform 1 0 88 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1683038052
transform 1 0 96 0 1 1570
box -8 -3 104 105
use M3_M2  M3_M2_51
timestamp 1683038052
transform 1 0 204 0 1 1575
box -3 -3 3 3
use FILL  FILL_3
timestamp 1683038052
transform 1 0 192 0 1 1570
box -8 -3 16 105
use FILL  FILL_4
timestamp 1683038052
transform 1 0 200 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_52
timestamp 1683038052
transform 1 0 236 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1683038052
transform 1 0 284 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_1
timestamp 1683038052
transform -1 0 304 0 1 1570
box -8 -3 104 105
use FILL  FILL_5
timestamp 1683038052
transform 1 0 304 0 1 1570
box -8 -3 16 105
use FILL  FILL_6
timestamp 1683038052
transform 1 0 312 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1683038052
transform 1 0 320 0 1 1570
box -8 -3 104 105
use FILL  FILL_7
timestamp 1683038052
transform 1 0 416 0 1 1570
box -8 -3 16 105
use FILL  FILL_8
timestamp 1683038052
transform 1 0 424 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_0
timestamp 1683038052
transform 1 0 432 0 1 1570
box -8 -3 40 105
use OAI21X1  OAI21X1_0
timestamp 1683038052
transform 1 0 464 0 1 1570
box -8 -3 34 105
use NAND3X1  NAND3X1_1
timestamp 1683038052
transform 1 0 496 0 1 1570
box -8 -3 40 105
use OAI21X1  OAI21X1_1
timestamp 1683038052
transform 1 0 528 0 1 1570
box -8 -3 34 105
use FILL  FILL_9
timestamp 1683038052
transform 1 0 560 0 1 1570
box -8 -3 16 105
use FILL  FILL_10
timestamp 1683038052
transform 1 0 568 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1683038052
transform 1 0 576 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1683038052
transform 1 0 672 0 1 1570
box -8 -3 104 105
use FILL  FILL_11
timestamp 1683038052
transform 1 0 768 0 1 1570
box -8 -3 16 105
use FILL  FILL_12
timestamp 1683038052
transform 1 0 776 0 1 1570
box -8 -3 16 105
use FILL  FILL_20
timestamp 1683038052
transform 1 0 784 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_6
timestamp 1683038052
transform 1 0 792 0 1 1570
box -9 -3 26 105
use NAND3X1  NAND3X1_5
timestamp 1683038052
transform 1 0 808 0 1 1570
box -8 -3 40 105
use FILL  FILL_22
timestamp 1683038052
transform 1 0 840 0 1 1570
box -8 -3 16 105
use FILL  FILL_23
timestamp 1683038052
transform 1 0 848 0 1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_6
timestamp 1683038052
transform 1 0 856 0 1 1570
box -8 -3 34 105
use NAND2X1  NAND2X1_3
timestamp 1683038052
transform 1 0 888 0 1 1570
box -8 -3 32 105
use FILL  FILL_25
timestamp 1683038052
transform 1 0 912 0 1 1570
box -8 -3 16 105
use FILL  FILL_31
timestamp 1683038052
transform 1 0 920 0 1 1570
box -8 -3 16 105
use FILL  FILL_32
timestamp 1683038052
transform 1 0 928 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_54
timestamp 1683038052
transform 1 0 964 0 1 1575
box -3 -3 3 3
use OAI21X1  OAI21X1_7
timestamp 1683038052
transform 1 0 936 0 1 1570
box -8 -3 34 105
use FILL  FILL_33
timestamp 1683038052
transform 1 0 968 0 1 1570
box -8 -3 16 105
use FAX1  FAX1_0
timestamp 1683038052
transform 1 0 976 0 1 1570
box -5 -3 126 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1683038052
transform -1 0 1192 0 1 1570
box -8 -3 104 105
use FILL  FILL_37
timestamp 1683038052
transform 1 0 1192 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_7
timestamp 1683038052
transform 1 0 1200 0 1 1570
box -9 -3 26 105
use FAX1  FAX1_1
timestamp 1683038052
transform 1 0 1216 0 1 1570
box -5 -3 126 105
use M3_M2  M3_M2_55
timestamp 1683038052
transform 1 0 1348 0 1 1575
box -3 -3 3 3
use INVX2  INVX2_8
timestamp 1683038052
transform -1 0 1352 0 1 1570
box -9 -3 26 105
use FILL  FILL_38
timestamp 1683038052
transform 1 0 1352 0 1 1570
box -8 -3 16 105
use FILL  FILL_39
timestamp 1683038052
transform 1 0 1360 0 1 1570
box -8 -3 16 105
use FILL  FILL_40
timestamp 1683038052
transform 1 0 1368 0 1 1570
box -8 -3 16 105
use FILL  FILL_41
timestamp 1683038052
transform 1 0 1376 0 1 1570
box -8 -3 16 105
use FAX1  FAX1_2
timestamp 1683038052
transform 1 0 1384 0 1 1570
box -5 -3 126 105
use FILL  FILL_42
timestamp 1683038052
transform 1 0 1504 0 1 1570
box -8 -3 16 105
use FILL  FILL_43
timestamp 1683038052
transform 1 0 1512 0 1 1570
box -8 -3 16 105
use FILL  FILL_66
timestamp 1683038052
transform 1 0 1520 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_12
timestamp 1683038052
transform 1 0 1528 0 1 1570
box -9 -3 26 105
use FILL  FILL_68
timestamp 1683038052
transform 1 0 1544 0 1 1570
box -8 -3 16 105
use FILL  FILL_72
timestamp 1683038052
transform 1 0 1552 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1683038052
transform 1 0 1560 0 1 1570
box -8 -3 104 105
use FILL  FILL_74
timestamp 1683038052
transform 1 0 1656 0 1 1570
box -8 -3 16 105
use FILL  FILL_84
timestamp 1683038052
transform 1 0 1664 0 1 1570
box -8 -3 16 105
use FILL  FILL_86
timestamp 1683038052
transform 1 0 1672 0 1 1570
box -8 -3 16 105
use FILL  FILL_88
timestamp 1683038052
transform 1 0 1680 0 1 1570
box -8 -3 16 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_3
timestamp 1683038052
transform 1 0 1716 0 1 1570
box -10 -3 10 3
use M2_M1  M2_M1_73
timestamp 1683038052
transform 1 0 76 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_77
timestamp 1683038052
transform 1 0 84 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1683038052
transform 1 0 108 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_74
timestamp 1683038052
transform 1 0 124 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1683038052
transform 1 0 84 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1683038052
transform 1 0 100 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_86
timestamp 1683038052
transform 1 0 124 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_75
timestamp 1683038052
transform 1 0 148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1683038052
transform 1 0 132 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1683038052
transform 1 0 148 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_150
timestamp 1683038052
transform 1 0 100 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1683038052
transform 1 0 116 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_120
timestamp 1683038052
transform 1 0 84 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_166
timestamp 1683038052
transform 1 0 92 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_100
timestamp 1683038052
transform 1 0 132 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_152
timestamp 1683038052
transform 1 0 148 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1683038052
transform 1 0 156 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_121
timestamp 1683038052
transform 1 0 156 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_113
timestamp 1683038052
transform 1 0 188 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1683038052
transform 1 0 180 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_101
timestamp 1683038052
transform 1 0 188 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_154
timestamp 1683038052
transform 1 0 196 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_122
timestamp 1683038052
transform 1 0 180 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_77
timestamp 1683038052
transform 1 0 212 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1683038052
transform 1 0 212 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_123
timestamp 1683038052
transform 1 0 212 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_78
timestamp 1683038052
transform 1 0 236 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1683038052
transform 1 0 260 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1683038052
transform 1 0 276 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1683038052
transform 1 0 284 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1683038052
transform 1 0 252 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1683038052
transform 1 0 260 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_87
timestamp 1683038052
transform 1 0 284 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_117
timestamp 1683038052
transform 1 0 292 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_124
timestamp 1683038052
transform 1 0 276 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_81
timestamp 1683038052
transform 1 0 324 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1683038052
transform 1 0 308 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_88
timestamp 1683038052
transform 1 0 332 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_119
timestamp 1683038052
transform 1 0 340 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_102
timestamp 1683038052
transform 1 0 308 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_155
timestamp 1683038052
transform 1 0 324 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_156
timestamp 1683038052
transform 1 0 332 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_103
timestamp 1683038052
transform 1 0 340 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1683038052
transform 1 0 364 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_82
timestamp 1683038052
transform 1 0 364 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1683038052
transform 1 0 356 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_125
timestamp 1683038052
transform 1 0 324 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_167
timestamp 1683038052
transform 1 0 348 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_126
timestamp 1683038052
transform 1 0 356 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1683038052
transform 1 0 380 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_57
timestamp 1683038052
transform 1 0 428 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_62
timestamp 1683038052
transform 1 0 420 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1683038052
transform 1 0 444 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_83
timestamp 1683038052
transform 1 0 428 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1683038052
transform 1 0 444 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1683038052
transform 1 0 460 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_79
timestamp 1683038052
transform 1 0 476 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_86
timestamp 1683038052
transform 1 0 484 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1683038052
transform 1 0 428 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1683038052
transform 1 0 436 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1683038052
transform 1 0 452 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_89
timestamp 1683038052
transform 1 0 460 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1683038052
transform 1 0 452 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1683038052
transform 1 0 428 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1683038052
transform 1 0 468 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_80
timestamp 1683038052
transform 1 0 500 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_87
timestamp 1683038052
transform 1 0 524 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_90
timestamp 1683038052
transform 1 0 492 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_123
timestamp 1683038052
transform 1 0 500 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1683038052
transform 1 0 492 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1683038052
transform 1 0 548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1683038052
transform 1 0 532 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1683038052
transform 1 0 548 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1683038052
transform 1 0 516 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_104
timestamp 1683038052
transform 1 0 524 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_168
timestamp 1683038052
transform 1 0 508 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1683038052
transform 1 0 548 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_128
timestamp 1683038052
transform 1 0 548 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1683038052
transform 1 0 532 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1683038052
transform 1 0 628 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_69
timestamp 1683038052
transform 1 0 668 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1683038052
transform 1 0 700 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_71
timestamp 1683038052
transform 1 0 732 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_89
timestamp 1683038052
transform 1 0 652 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_81
timestamp 1683038052
transform 1 0 668 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1683038052
transform 1 0 772 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_90
timestamp 1683038052
transform 1 0 748 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1683038052
transform 1 0 764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1683038052
transform 1 0 564 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1683038052
transform 1 0 628 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_91
timestamp 1683038052
transform 1 0 652 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_128
timestamp 1683038052
transform 1 0 668 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_105
timestamp 1683038052
transform 1 0 564 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1683038052
transform 1 0 652 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1683038052
transform 1 0 684 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_129
timestamp 1683038052
transform 1 0 724 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_93
timestamp 1683038052
transform 1 0 748 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1683038052
transform 1 0 676 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1683038052
transform 1 0 724 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1683038052
transform 1 0 764 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1683038052
transform 1 0 764 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_92
timestamp 1683038052
transform 1 0 780 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_82
timestamp 1683038052
transform 1 0 788 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_130
timestamp 1683038052
transform 1 0 788 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_73
timestamp 1683038052
transform 1 0 820 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_93
timestamp 1683038052
transform 1 0 820 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_94
timestamp 1683038052
transform 1 0 812 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_131
timestamp 1683038052
transform 1 0 820 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1683038052
transform 1 0 828 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1683038052
transform 1 0 812 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_110
timestamp 1683038052
transform 1 0 836 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_94
timestamp 1683038052
transform 1 0 860 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_95
timestamp 1683038052
transform 1 0 852 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_162
timestamp 1683038052
transform 1 0 844 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1683038052
transform 1 0 852 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_83
timestamp 1683038052
transform 1 0 876 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_95
timestamp 1683038052
transform 1 0 884 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1683038052
transform 1 0 868 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_96
timestamp 1683038052
transform 1 0 876 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1683038052
transform 1 0 900 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_134
timestamp 1683038052
transform 1 0 892 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_111
timestamp 1683038052
transform 1 0 892 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_96
timestamp 1683038052
transform 1 0 908 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_130
timestamp 1683038052
transform 1 0 908 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_63
timestamp 1683038052
transform 1 0 948 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_164
timestamp 1683038052
transform 1 0 948 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1683038052
transform 1 0 988 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1683038052
transform 1 0 1004 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1683038052
transform 1 0 1020 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_84
timestamp 1683038052
transform 1 0 1084 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_99
timestamp 1683038052
transform 1 0 1124 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1683038052
transform 1 0 1140 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_85
timestamp 1683038052
transform 1 0 1148 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_136
timestamp 1683038052
transform 1 0 1108 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1683038052
transform 1 0 1116 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1683038052
transform 1 0 1132 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1683038052
transform 1 0 1148 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_112
timestamp 1683038052
transform 1 0 1108 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_131
timestamp 1683038052
transform 1 0 1124 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1683038052
transform 1 0 1140 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1683038052
transform 1 0 1284 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_59
timestamp 1683038052
transform 1 0 1356 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_64
timestamp 1683038052
transform 1 0 1172 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_65
timestamp 1683038052
transform 1 0 1196 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_75
timestamp 1683038052
transform 1 0 1164 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_76
timestamp 1683038052
transform 1 0 1220 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_71
timestamp 1683038052
transform 1 0 1268 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1683038052
transform 1 0 1388 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1683038052
transform 1 0 1164 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1683038052
transform 1 0 1276 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1683038052
transform 1 0 1284 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1683038052
transform 1 0 1172 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1683038052
transform 1 0 1180 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_97
timestamp 1683038052
transform 1 0 1268 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1683038052
transform 1 0 1284 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_142
timestamp 1683038052
transform 1 0 1292 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_143
timestamp 1683038052
transform 1 0 1300 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_99
timestamp 1683038052
transform 1 0 1324 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_113
timestamp 1683038052
transform 1 0 1172 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_114
timestamp 1683038052
transform 1 0 1276 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_115
timestamp 1683038052
transform 1 0 1300 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_132
timestamp 1683038052
transform 1 0 1188 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1683038052
transform 1 0 1252 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1683038052
transform 1 0 1276 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_144
timestamp 1683038052
transform 1 0 1404 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1683038052
transform 1 0 1412 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1683038052
transform 1 0 1428 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1683038052
transform 1 0 1452 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_145
timestamp 1683038052
transform 1 0 1444 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_116
timestamp 1683038052
transform 1 0 1444 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1683038052
transform 1 0 1452 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_146
timestamp 1683038052
transform 1 0 1484 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1683038052
transform 1 0 1492 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_117
timestamp 1683038052
transform 1 0 1492 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1683038052
transform 1 0 1532 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_147
timestamp 1683038052
transform 1 0 1524 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_118
timestamp 1683038052
transform 1 0 1556 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_165
timestamp 1683038052
transform 1 0 1564 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1683038052
transform 1 0 1580 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1683038052
transform 1 0 1596 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_119
timestamp 1683038052
transform 1 0 1596 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_149
timestamp 1683038052
transform 1 0 1636 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_61
timestamp 1683038052
transform 1 0 1652 0 1 1565
box -3 -3 3 3
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_4
timestamp 1683038052
transform 1 0 24 0 1 1470
box -10 -3 10 3
use INVX2  INVX2_0
timestamp 1683038052
transform 1 0 72 0 -1 1570
box -9 -3 26 105
use NAND3X1  NAND3X1_2
timestamp 1683038052
transform 1 0 88 0 -1 1570
box -8 -3 40 105
use OAI21X1  OAI21X1_2
timestamp 1683038052
transform 1 0 120 0 -1 1570
box -8 -3 34 105
use FILL  FILL_13
timestamp 1683038052
transform 1 0 152 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_0
timestamp 1683038052
transform 1 0 160 0 -1 1570
box -8 -3 32 105
use FILL  FILL_14
timestamp 1683038052
transform 1 0 184 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_1
timestamp 1683038052
transform -1 0 216 0 -1 1570
box -8 -3 32 105
use INVX2  INVX2_1
timestamp 1683038052
transform 1 0 216 0 -1 1570
box -9 -3 26 105
use FILL  FILL_15
timestamp 1683038052
transform 1 0 232 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_2
timestamp 1683038052
transform 1 0 240 0 -1 1570
box -9 -3 26 105
use AOI21X1  AOI21X1_0
timestamp 1683038052
transform -1 0 288 0 -1 1570
box -7 -3 39 105
use FILL  FILL_16
timestamp 1683038052
transform 1 0 288 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_3
timestamp 1683038052
transform 1 0 296 0 -1 1570
box -8 -3 34 105
use NAND3X1  NAND3X1_3
timestamp 1683038052
transform 1 0 328 0 -1 1570
box -8 -3 40 105
use FILL  FILL_17
timestamp 1683038052
transform 1 0 360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_18
timestamp 1683038052
transform 1 0 368 0 -1 1570
box -8 -3 16 105
use XOR2X1  XOR2X1_0
timestamp 1683038052
transform 1 0 376 0 -1 1570
box -8 -3 64 105
use AOI22X1  AOI22X1_0
timestamp 1683038052
transform 1 0 432 0 -1 1570
box -8 -3 46 105
use INVX2  INVX2_3
timestamp 1683038052
transform -1 0 488 0 -1 1570
box -9 -3 26 105
use NAND3X1  NAND3X1_4
timestamp 1683038052
transform 1 0 488 0 -1 1570
box -8 -3 40 105
use OAI21X1  OAI21X1_4
timestamp 1683038052
transform 1 0 520 0 -1 1570
box -8 -3 34 105
use INVX2  INVX2_4
timestamp 1683038052
transform -1 0 568 0 -1 1570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1683038052
transform -1 0 664 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1683038052
transform -1 0 760 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_5
timestamp 1683038052
transform 1 0 760 0 -1 1570
box -9 -3 26 105
use FILL  FILL_19
timestamp 1683038052
transform 1 0 776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_21
timestamp 1683038052
transform 1 0 784 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_2
timestamp 1683038052
transform 1 0 792 0 -1 1570
box -8 -3 32 105
use OAI21X1  OAI21X1_5
timestamp 1683038052
transform 1 0 816 0 -1 1570
box -8 -3 34 105
use FILL  FILL_24
timestamp 1683038052
transform 1 0 848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_26
timestamp 1683038052
transform 1 0 856 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_4
timestamp 1683038052
transform -1 0 888 0 -1 1570
box -8 -3 32 105
use FILL  FILL_27
timestamp 1683038052
transform 1 0 888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_28
timestamp 1683038052
transform 1 0 896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_29
timestamp 1683038052
transform 1 0 904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_30
timestamp 1683038052
transform 1 0 912 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_8
timestamp 1683038052
transform 1 0 920 0 -1 1570
box -8 -3 34 105
use FILL  FILL_34
timestamp 1683038052
transform 1 0 952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_35
timestamp 1683038052
transform 1 0 960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_36
timestamp 1683038052
transform 1 0 968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_44
timestamp 1683038052
transform 1 0 976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_45
timestamp 1683038052
transform 1 0 984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_46
timestamp 1683038052
transform 1 0 992 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_9
timestamp 1683038052
transform 1 0 1000 0 -1 1570
box -9 -3 26 105
use FILL  FILL_47
timestamp 1683038052
transform 1 0 1016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_48
timestamp 1683038052
transform 1 0 1024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_49
timestamp 1683038052
transform 1 0 1032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_50
timestamp 1683038052
transform 1 0 1040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_51
timestamp 1683038052
transform 1 0 1048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_52
timestamp 1683038052
transform 1 0 1056 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_10
timestamp 1683038052
transform 1 0 1064 0 -1 1570
box -9 -3 26 105
use FILL  FILL_53
timestamp 1683038052
transform 1 0 1080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_54
timestamp 1683038052
transform 1 0 1088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_55
timestamp 1683038052
transform 1 0 1096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_56
timestamp 1683038052
transform 1 0 1104 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_1
timestamp 1683038052
transform -1 0 1152 0 -1 1570
box -8 -3 46 105
use FILL  FILL_57
timestamp 1683038052
transform 1 0 1152 0 -1 1570
box -8 -3 16 105
use FAX1  FAX1_3
timestamp 1683038052
transform 1 0 1160 0 -1 1570
box -5 -3 126 105
use FAX1  FAX1_4
timestamp 1683038052
transform 1 0 1280 0 -1 1570
box -5 -3 126 105
use FILL  FILL_58
timestamp 1683038052
transform 1 0 1400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_59
timestamp 1683038052
transform 1 0 1408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_60
timestamp 1683038052
transform 1 0 1416 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_2
timestamp 1683038052
transform -1 0 1464 0 -1 1570
box -8 -3 46 105
use FILL  FILL_61
timestamp 1683038052
transform 1 0 1464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_62
timestamp 1683038052
transform 1 0 1472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_63
timestamp 1683038052
transform 1 0 1480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_64
timestamp 1683038052
transform 1 0 1488 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_11
timestamp 1683038052
transform 1 0 1496 0 -1 1570
box -9 -3 26 105
use FILL  FILL_65
timestamp 1683038052
transform 1 0 1512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_67
timestamp 1683038052
transform 1 0 1520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_69
timestamp 1683038052
transform 1 0 1528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_70
timestamp 1683038052
transform 1 0 1536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_71
timestamp 1683038052
transform 1 0 1544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_73
timestamp 1683038052
transform 1 0 1552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_75
timestamp 1683038052
transform 1 0 1560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_76
timestamp 1683038052
transform 1 0 1568 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_9
timestamp 1683038052
transform -1 0 1608 0 -1 1570
box -8 -3 34 105
use FILL  FILL_77
timestamp 1683038052
transform 1 0 1608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_78
timestamp 1683038052
transform 1 0 1616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_79
timestamp 1683038052
transform 1 0 1624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_80
timestamp 1683038052
transform 1 0 1632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_81
timestamp 1683038052
transform 1 0 1640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_82
timestamp 1683038052
transform 1 0 1648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_83
timestamp 1683038052
transform 1 0 1656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_85
timestamp 1683038052
transform 1 0 1664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_87
timestamp 1683038052
transform 1 0 1672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_89
timestamp 1683038052
transform 1 0 1680 0 -1 1570
box -8 -3 16 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_5
timestamp 1683038052
transform 1 0 1740 0 1 1470
box -10 -3 10 3
use M2_M1  M2_M1_185
timestamp 1683038052
transform 1 0 76 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_150
timestamp 1683038052
transform 1 0 108 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1683038052
transform 1 0 132 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_186
timestamp 1683038052
transform 1 0 132 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_143
timestamp 1683038052
transform 1 0 156 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_169
timestamp 1683038052
transform 1 0 156 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1683038052
transform 1 0 148 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1683038052
transform 1 0 140 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_178
timestamp 1683038052
transform 1 0 140 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1683038052
transform 1 0 164 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1683038052
transform 1 0 196 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_170
timestamp 1683038052
transform 1 0 188 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1683038052
transform 1 0 172 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_175
timestamp 1683038052
transform 1 0 180 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_158
timestamp 1683038052
transform 1 0 188 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_176
timestamp 1683038052
transform 1 0 196 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1683038052
transform 1 0 164 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_165
timestamp 1683038052
transform 1 0 172 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_188
timestamp 1683038052
transform 1 0 196 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_179
timestamp 1683038052
transform 1 0 164 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1683038052
transform 1 0 204 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_189
timestamp 1683038052
transform 1 0 212 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_151
timestamp 1683038052
transform 1 0 332 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_159
timestamp 1683038052
transform 1 0 340 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1683038052
transform 1 0 380 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_190
timestamp 1683038052
transform 1 0 268 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1683038052
transform 1 0 332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1683038052
transform 1 0 340 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1683038052
transform 1 0 380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1683038052
transform 1 0 444 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1683038052
transform 1 0 316 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_186
timestamp 1683038052
transform 1 0 324 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_226
timestamp 1683038052
transform 1 0 428 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1683038052
transform 1 0 444 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_187
timestamp 1683038052
transform 1 0 380 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1683038052
transform 1 0 428 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1683038052
transform 1 0 452 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_195
timestamp 1683038052
transform 1 0 460 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1683038052
transform 1 0 460 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1683038052
transform 1 0 492 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_174
timestamp 1683038052
transform 1 0 492 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_197
timestamp 1683038052
transform 1 0 508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1683038052
transform 1 0 516 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1683038052
transform 1 0 508 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_175
timestamp 1683038052
transform 1 0 516 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_199
timestamp 1683038052
transform 1 0 540 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1683038052
transform 1 0 524 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1683038052
transform 1 0 548 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_141
timestamp 1683038052
transform 1 0 564 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_177
timestamp 1683038052
transform 1 0 564 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1683038052
transform 1 0 556 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_144
timestamp 1683038052
transform 1 0 604 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_171
timestamp 1683038052
transform 1 0 612 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_178
timestamp 1683038052
transform 1 0 612 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1683038052
transform 1 0 604 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_167
timestamp 1683038052
transform 1 0 612 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_232
timestamp 1683038052
transform 1 0 620 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1683038052
transform 1 0 620 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1683038052
transform 1 0 636 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1683038052
transform 1 0 676 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_168
timestamp 1683038052
transform 1 0 724 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1683038052
transform 1 0 748 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_204
timestamp 1683038052
transform 1 0 732 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1683038052
transform 1 0 652 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_189
timestamp 1683038052
transform 1 0 644 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1683038052
transform 1 0 684 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1683038052
transform 1 0 756 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_205
timestamp 1683038052
transform 1 0 764 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1683038052
transform 1 0 748 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1683038052
transform 1 0 756 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_145
timestamp 1683038052
transform 1 0 788 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_172
timestamp 1683038052
transform 1 0 780 0 1 1435
box -2 -2 2 2
use M3_M2  M3_M2_163
timestamp 1683038052
transform 1 0 780 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1683038052
transform 1 0 796 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_179
timestamp 1683038052
transform 1 0 788 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1683038052
transform 1 0 804 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1683038052
transform 1 0 796 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1683038052
transform 1 0 812 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1683038052
transform 1 0 836 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_146
timestamp 1683038052
transform 1 0 852 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_181
timestamp 1683038052
transform 1 0 852 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_153
timestamp 1683038052
transform 1 0 868 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_182
timestamp 1683038052
transform 1 0 868 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_170
timestamp 1683038052
transform 1 0 860 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_237
timestamp 1683038052
transform 1 0 876 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_171
timestamp 1683038052
transform 1 0 908 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_238
timestamp 1683038052
transform 1 0 900 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1683038052
transform 1 0 908 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_154
timestamp 1683038052
transform 1 0 932 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1683038052
transform 1 0 956 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_183
timestamp 1683038052
transform 1 0 932 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_164
timestamp 1683038052
transform 1 0 940 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_208
timestamp 1683038052
transform 1 0 940 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1683038052
transform 1 0 956 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1683038052
transform 1 0 972 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1683038052
transform 1 0 964 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_155
timestamp 1683038052
transform 1 0 1004 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_211
timestamp 1683038052
transform 1 0 1004 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_180
timestamp 1683038052
transform 1 0 996 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_212
timestamp 1683038052
transform 1 0 1028 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1683038052
transform 1 0 1012 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_181
timestamp 1683038052
transform 1 0 1092 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_253
timestamp 1683038052
transform 1 0 1116 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1683038052
transform 1 0 1140 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_172
timestamp 1683038052
transform 1 0 1148 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_242
timestamp 1683038052
transform 1 0 1148 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_148
timestamp 1683038052
transform 1 0 1164 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_213
timestamp 1683038052
transform 1 0 1172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1683038052
transform 1 0 1156 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_173
timestamp 1683038052
transform 1 0 1180 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1683038052
transform 1 0 1196 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_244
timestamp 1683038052
transform 1 0 1180 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1683038052
transform 1 0 1188 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_182
timestamp 1683038052
transform 1 0 1180 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1683038052
transform 1 0 1204 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_214
timestamp 1683038052
transform 1 0 1252 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1683038052
transform 1 0 1268 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1683038052
transform 1 0 1284 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1683038052
transform 1 0 1260 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1683038052
transform 1 0 1276 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_191
timestamp 1683038052
transform 1 0 1260 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1683038052
transform 1 0 1420 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_217
timestamp 1683038052
transform 1 0 1412 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1683038052
transform 1 0 1420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1683038052
transform 1 0 1316 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1683038052
transform 1 0 1324 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_192
timestamp 1683038052
transform 1 0 1332 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1683038052
transform 1 0 1356 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1683038052
transform 1 0 1420 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_249
timestamp 1683038052
transform 1 0 1436 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_195
timestamp 1683038052
transform 1 0 1436 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_219
timestamp 1683038052
transform 1 0 1484 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_176
timestamp 1683038052
transform 1 0 1484 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_220
timestamp 1683038052
transform 1 0 1524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1683038052
transform 1 0 1580 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1683038052
transform 1 0 1500 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_177
timestamp 1683038052
transform 1 0 1524 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1683038052
transform 1 0 1516 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1683038052
transform 1 0 1532 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1683038052
transform 1 0 1532 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_222
timestamp 1683038052
transform 1 0 1628 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1683038052
transform 1 0 1692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1683038052
transform 1 0 1604 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_197
timestamp 1683038052
transform 1 0 1644 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1683038052
transform 1 0 1692 0 1 1385
box -3 -3 3 3
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_6
timestamp 1683038052
transform 1 0 48 0 1 1370
box -10 -3 10 3
use FILL  FILL_90
timestamp 1683038052
transform 1 0 72 0 1 1370
box -8 -3 16 105
use FILL  FILL_92
timestamp 1683038052
transform 1 0 80 0 1 1370
box -8 -3 16 105
use FILL  FILL_93
timestamp 1683038052
transform 1 0 88 0 1 1370
box -8 -3 16 105
use FILL  FILL_94
timestamp 1683038052
transform 1 0 96 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_13
timestamp 1683038052
transform -1 0 120 0 1 1370
box -9 -3 26 105
use FILL  FILL_95
timestamp 1683038052
transform 1 0 120 0 1 1370
box -8 -3 16 105
use FILL  FILL_96
timestamp 1683038052
transform 1 0 128 0 1 1370
box -8 -3 16 105
use FILL  FILL_97
timestamp 1683038052
transform 1 0 136 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_6
timestamp 1683038052
transform -1 0 176 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_7
timestamp 1683038052
transform -1 0 208 0 1 1370
box -8 -3 40 105
use FILL  FILL_98
timestamp 1683038052
transform 1 0 208 0 1 1370
box -8 -3 16 105
use FILL  FILL_103
timestamp 1683038052
transform 1 0 216 0 1 1370
box -8 -3 16 105
use FILL  FILL_105
timestamp 1683038052
transform 1 0 224 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1683038052
transform -1 0 328 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_15
timestamp 1683038052
transform -1 0 344 0 1 1370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1683038052
transform -1 0 440 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_16
timestamp 1683038052
transform 1 0 440 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_17
timestamp 1683038052
transform 1 0 456 0 1 1370
box -9 -3 26 105
use FILL  FILL_106
timestamp 1683038052
transform 1 0 472 0 1 1370
box -8 -3 16 105
use FILL  FILL_115
timestamp 1683038052
transform 1 0 480 0 1 1370
box -8 -3 16 105
use FILL  FILL_117
timestamp 1683038052
transform 1 0 488 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_20
timestamp 1683038052
transform -1 0 512 0 1 1370
box -9 -3 26 105
use AOI21X1  AOI21X1_2
timestamp 1683038052
transform 1 0 512 0 1 1370
box -7 -3 39 105
use INVX2  INVX2_21
timestamp 1683038052
transform 1 0 544 0 1 1370
box -9 -3 26 105
use FILL  FILL_118
timestamp 1683038052
transform 1 0 560 0 1 1370
box -8 -3 16 105
use FILL  FILL_119
timestamp 1683038052
transform 1 0 568 0 1 1370
box -8 -3 16 105
use FILL  FILL_120
timestamp 1683038052
transform 1 0 576 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_8
timestamp 1683038052
transform -1 0 616 0 1 1370
box -8 -3 40 105
use NOR2X1  NOR2X1_0
timestamp 1683038052
transform 1 0 616 0 1 1370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1683038052
transform 1 0 640 0 1 1370
box -8 -3 104 105
use NOR2X1  NOR2X1_1
timestamp 1683038052
transform 1 0 736 0 1 1370
box -8 -3 32 105
use INVX2  INVX2_22
timestamp 1683038052
transform 1 0 760 0 1 1370
box -9 -3 26 105
use FILL  FILL_124
timestamp 1683038052
transform 1 0 776 0 1 1370
box -8 -3 16 105
use FILL  FILL_125
timestamp 1683038052
transform 1 0 784 0 1 1370
box -8 -3 16 105
use FILL  FILL_126
timestamp 1683038052
transform 1 0 792 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_9
timestamp 1683038052
transform 1 0 800 0 1 1370
box -8 -3 40 105
use FILL  FILL_127
timestamp 1683038052
transform 1 0 832 0 1 1370
box -8 -3 16 105
use FILL  FILL_133
timestamp 1683038052
transform 1 0 840 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_9
timestamp 1683038052
transform 1 0 848 0 1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_12
timestamp 1683038052
transform 1 0 872 0 1 1370
box -8 -3 34 105
use FILL  FILL_135
timestamp 1683038052
transform 1 0 904 0 1 1370
box -8 -3 16 105
use FILL  FILL_141
timestamp 1683038052
transform 1 0 912 0 1 1370
box -8 -3 16 105
use FILL  FILL_142
timestamp 1683038052
transform 1 0 920 0 1 1370
box -8 -3 16 105
use AND2X2  AND2X2_0
timestamp 1683038052
transform 1 0 928 0 1 1370
box -8 -3 40 105
use FILL  FILL_143
timestamp 1683038052
transform 1 0 960 0 1 1370
box -8 -3 16 105
use FILL  FILL_144
timestamp 1683038052
transform 1 0 968 0 1 1370
box -8 -3 16 105
use FILL  FILL_145
timestamp 1683038052
transform 1 0 976 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_25
timestamp 1683038052
transform 1 0 984 0 1 1370
box -9 -3 26 105
use FILL  FILL_146
timestamp 1683038052
transform 1 0 1000 0 1 1370
box -8 -3 16 105
use FAX1  FAX1_5
timestamp 1683038052
transform 1 0 1008 0 1 1370
box -5 -3 126 105
use FILL  FILL_147
timestamp 1683038052
transform 1 0 1128 0 1 1370
box -8 -3 16 105
use FILL  FILL_148
timestamp 1683038052
transform 1 0 1136 0 1 1370
box -8 -3 16 105
use FILL  FILL_149
timestamp 1683038052
transform 1 0 1144 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_13
timestamp 1683038052
transform -1 0 1184 0 1 1370
box -8 -3 34 105
use FILL  FILL_150
timestamp 1683038052
transform 1 0 1184 0 1 1370
box -8 -3 16 105
use FILL  FILL_151
timestamp 1683038052
transform 1 0 1192 0 1 1370
box -8 -3 16 105
use FILL  FILL_155
timestamp 1683038052
transform 1 0 1200 0 1 1370
box -8 -3 16 105
use FILL  FILL_157
timestamp 1683038052
transform 1 0 1208 0 1 1370
box -8 -3 16 105
use FILL  FILL_158
timestamp 1683038052
transform 1 0 1216 0 1 1370
box -8 -3 16 105
use FILL  FILL_159
timestamp 1683038052
transform 1 0 1224 0 1 1370
box -8 -3 16 105
use FILL  FILL_160
timestamp 1683038052
transform 1 0 1232 0 1 1370
box -8 -3 16 105
use FILL  FILL_161
timestamp 1683038052
transform 1 0 1240 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_3
timestamp 1683038052
transform -1 0 1288 0 1 1370
box -8 -3 46 105
use FILL  FILL_162
timestamp 1683038052
transform 1 0 1288 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_199
timestamp 1683038052
transform 1 0 1308 0 1 1375
box -3 -3 3 3
use FILL  FILL_163
timestamp 1683038052
transform 1 0 1296 0 1 1370
box -8 -3 16 105
use FILL  FILL_164
timestamp 1683038052
transform 1 0 1304 0 1 1370
box -8 -3 16 105
use FAX1  FAX1_7
timestamp 1683038052
transform -1 0 1432 0 1 1370
box -5 -3 126 105
use FILL  FILL_165
timestamp 1683038052
transform 1 0 1432 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_27
timestamp 1683038052
transform 1 0 1440 0 1 1370
box -9 -3 26 105
use FILL  FILL_166
timestamp 1683038052
transform 1 0 1456 0 1 1370
box -8 -3 16 105
use FILL  FILL_167
timestamp 1683038052
transform 1 0 1464 0 1 1370
box -8 -3 16 105
use FILL  FILL_168
timestamp 1683038052
transform 1 0 1472 0 1 1370
box -8 -3 16 105
use FILL  FILL_169
timestamp 1683038052
transform 1 0 1480 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_200
timestamp 1683038052
transform 1 0 1572 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_15
timestamp 1683038052
transform 1 0 1488 0 1 1370
box -8 -3 104 105
use FILL  FILL_170
timestamp 1683038052
transform 1 0 1584 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_201
timestamp 1683038052
transform 1 0 1604 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_17
timestamp 1683038052
transform 1 0 1592 0 1 1370
box -8 -3 104 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_7
timestamp 1683038052
transform 1 0 1716 0 1 1370
box -10 -3 10 3
use M2_M1  M2_M1_259
timestamp 1683038052
transform 1 0 84 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_225
timestamp 1683038052
transform 1 0 92 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_260
timestamp 1683038052
transform 1 0 108 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1683038052
transform 1 0 92 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1683038052
transform 1 0 116 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1683038052
transform 1 0 100 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_240
timestamp 1683038052
transform 1 0 116 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1683038052
transform 1 0 148 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_255
timestamp 1683038052
transform 1 0 164 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1683038052
transform 1 0 148 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1683038052
transform 1 0 132 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_250
timestamp 1683038052
transform 1 0 100 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_251
timestamp 1683038052
transform 1 0 132 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_262
timestamp 1683038052
transform 1 0 172 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1683038052
transform 1 0 164 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_209
timestamp 1683038052
transform 1 0 180 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1683038052
transform 1 0 180 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_300
timestamp 1683038052
transform 1 0 180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1683038052
transform 1 0 188 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_227
timestamp 1683038052
transform 1 0 196 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_241
timestamp 1683038052
transform 1 0 188 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_301
timestamp 1683038052
transform 1 0 228 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_204
timestamp 1683038052
transform 1 0 252 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_210
timestamp 1683038052
transform 1 0 276 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_264
timestamp 1683038052
transform 1 0 244 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_228
timestamp 1683038052
transform 1 0 252 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_265
timestamp 1683038052
transform 1 0 260 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1683038052
transform 1 0 276 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1683038052
transform 1 0 236 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_235
timestamp 1683038052
transform 1 0 244 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_303
timestamp 1683038052
transform 1 0 252 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1683038052
transform 1 0 268 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_252
timestamp 1683038052
transform 1 0 236 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_266
timestamp 1683038052
transform 1 0 268 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1683038052
transform 1 0 308 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1683038052
transform 1 0 300 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_267
timestamp 1683038052
transform 1 0 300 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1683038052
transform 1 0 324 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1683038052
transform 1 0 340 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1683038052
transform 1 0 292 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_242
timestamp 1683038052
transform 1 0 292 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_306
timestamp 1683038052
transform 1 0 332 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_236
timestamp 1683038052
transform 1 0 340 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_337
timestamp 1683038052
transform 1 0 300 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_243
timestamp 1683038052
transform 1 0 324 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_253
timestamp 1683038052
transform 1 0 300 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1683038052
transform 1 0 292 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_263
timestamp 1683038052
transform 1 0 308 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1683038052
transform 1 0 356 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_307
timestamp 1683038052
transform 1 0 356 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1683038052
transform 1 0 420 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1683038052
transform 1 0 396 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1683038052
transform 1 0 404 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_254
timestamp 1683038052
transform 1 0 396 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_271
timestamp 1683038052
transform 1 0 444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1683038052
transform 1 0 428 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_255
timestamp 1683038052
transform 1 0 428 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_267
timestamp 1683038052
transform 1 0 404 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_272
timestamp 1683038052
transform 1 0 492 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_229
timestamp 1683038052
transform 1 0 500 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_273
timestamp 1683038052
transform 1 0 508 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_230
timestamp 1683038052
transform 1 0 516 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_274
timestamp 1683038052
transform 1 0 524 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1683038052
transform 1 0 500 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1683038052
transform 1 0 516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1683038052
transform 1 0 532 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_244
timestamp 1683038052
transform 1 0 524 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_256
timestamp 1683038052
transform 1 0 516 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_275
timestamp 1683038052
transform 1 0 556 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1683038052
transform 1 0 556 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_257
timestamp 1683038052
transform 1 0 556 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1683038052
transform 1 0 596 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1683038052
transform 1 0 620 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_276
timestamp 1683038052
transform 1 0 644 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1683038052
transform 1 0 620 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_203
timestamp 1683038052
transform 1 0 676 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_277
timestamp 1683038052
transform 1 0 668 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1683038052
transform 1 0 692 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_245
timestamp 1683038052
transform 1 0 692 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1683038052
transform 1 0 756 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_278
timestamp 1683038052
transform 1 0 756 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_215
timestamp 1683038052
transform 1 0 780 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_279
timestamp 1683038052
transform 1 0 780 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1683038052
transform 1 0 780 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1683038052
transform 1 0 796 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1683038052
transform 1 0 820 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_216
timestamp 1683038052
transform 1 0 876 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_280
timestamp 1683038052
transform 1 0 876 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1683038052
transform 1 0 876 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1683038052
transform 1 0 884 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1683038052
transform 1 0 900 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1683038052
transform 1 0 924 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_231
timestamp 1683038052
transform 1 0 948 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_217
timestamp 1683038052
transform 1 0 956 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_281
timestamp 1683038052
transform 1 0 956 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_232
timestamp 1683038052
transform 1 0 964 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1683038052
transform 1 0 988 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_257
timestamp 1683038052
transform 1 0 1084 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1683038052
transform 1 0 980 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_233
timestamp 1683038052
transform 1 0 1084 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1683038052
transform 1 0 1180 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_283
timestamp 1683038052
transform 1 0 1092 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_234
timestamp 1683038052
transform 1 0 1108 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_284
timestamp 1683038052
transform 1 0 1180 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1683038052
transform 1 0 964 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1683038052
transform 1 0 972 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_323
timestamp 1683038052
transform 1 0 988 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_324
timestamp 1683038052
transform 1 0 996 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_246
timestamp 1683038052
transform 1 0 964 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1683038052
transform 1 0 1028 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1683038052
transform 1 0 1092 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_325
timestamp 1683038052
transform 1 0 1100 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1683038052
transform 1 0 1132 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_247
timestamp 1683038052
transform 1 0 996 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_258
timestamp 1683038052
transform 1 0 980 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_259
timestamp 1683038052
transform 1 0 1100 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1683038052
transform 1 0 1156 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_264
timestamp 1683038052
transform 1 0 1100 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_265
timestamp 1683038052
transform 1 0 1140 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1683038052
transform 1 0 1148 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_269
timestamp 1683038052
transform 1 0 1172 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_285
timestamp 1683038052
transform 1 0 1196 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1683038052
transform 1 0 1212 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_206
timestamp 1683038052
transform 1 0 1316 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1683038052
transform 1 0 1308 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_287
timestamp 1683038052
transform 1 0 1308 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1683038052
transform 1 0 1220 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1683038052
transform 1 0 1228 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1683038052
transform 1 0 1260 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_248
timestamp 1683038052
transform 1 0 1228 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_249
timestamp 1683038052
transform 1 0 1276 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_288
timestamp 1683038052
transform 1 0 1324 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_207
timestamp 1683038052
transform 1 0 1348 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1683038052
transform 1 0 1364 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_289
timestamp 1683038052
transform 1 0 1356 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1683038052
transform 1 0 1372 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1683038052
transform 1 0 1364 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1683038052
transform 1 0 1388 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1683038052
transform 1 0 1412 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1683038052
transform 1 0 1428 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_222
timestamp 1683038052
transform 1 0 1540 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_292
timestamp 1683038052
transform 1 0 1532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1683038052
transform 1 0 1540 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_239
timestamp 1683038052
transform 1 0 1500 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_332
timestamp 1683038052
transform 1 0 1516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1683038052
transform 1 0 1524 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1683038052
transform 1 0 1540 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_261
timestamp 1683038052
transform 1 0 1508 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_340
timestamp 1683038052
transform 1 0 1580 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_223
timestamp 1683038052
transform 1 0 1604 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_294
timestamp 1683038052
transform 1 0 1604 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_224
timestamp 1683038052
transform 1 0 1628 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_295
timestamp 1683038052
transform 1 0 1628 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1683038052
transform 1 0 1644 0 1 1335
box -2 -2 2 2
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_8
timestamp 1683038052
transform 1 0 24 0 1 1270
box -10 -3 10 3
use FILL  FILL_91
timestamp 1683038052
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_5
timestamp 1683038052
transform 1 0 80 0 -1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_10
timestamp 1683038052
transform 1 0 104 0 -1 1370
box -8 -3 34 105
use AOI21X1  AOI21X1_1
timestamp 1683038052
transform 1 0 136 0 -1 1370
box -7 -3 39 105
use FILL  FILL_99
timestamp 1683038052
transform 1 0 168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_100
timestamp 1683038052
transform 1 0 176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_101
timestamp 1683038052
transform 1 0 184 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_14
timestamp 1683038052
transform 1 0 192 0 -1 1370
box -9 -3 26 105
use FILL  FILL_102
timestamp 1683038052
transform 1 0 208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_104
timestamp 1683038052
transform 1 0 216 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_18
timestamp 1683038052
transform 1 0 224 0 -1 1370
box -9 -3 26 105
use OAI22X1  OAI22X1_0
timestamp 1683038052
transform -1 0 280 0 -1 1370
box -8 -3 46 105
use NAND2X1  NAND2X1_6
timestamp 1683038052
transform 1 0 280 0 -1 1370
box -8 -3 32 105
use OAI22X1  OAI22X1_1
timestamp 1683038052
transform 1 0 304 0 -1 1370
box -8 -3 46 105
use INVX2  INVX2_19
timestamp 1683038052
transform 1 0 344 0 -1 1370
box -9 -3 26 105
use FILL  FILL_107
timestamp 1683038052
transform 1 0 360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_108
timestamp 1683038052
transform 1 0 368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_109
timestamp 1683038052
transform 1 0 376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_110
timestamp 1683038052
transform 1 0 384 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_11
timestamp 1683038052
transform 1 0 392 0 -1 1370
box -8 -3 34 105
use NAND2X1  NAND2X1_7
timestamp 1683038052
transform -1 0 448 0 -1 1370
box -8 -3 32 105
use FILL  FILL_111
timestamp 1683038052
transform 1 0 448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_112
timestamp 1683038052
transform 1 0 456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_113
timestamp 1683038052
transform 1 0 464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_114
timestamp 1683038052
transform 1 0 472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_116
timestamp 1683038052
transform 1 0 480 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_23
timestamp 1683038052
transform 1 0 488 0 -1 1370
box -9 -3 26 105
use OAI22X1  OAI22X1_2
timestamp 1683038052
transform -1 0 544 0 -1 1370
box -8 -3 46 105
use FILL  FILL_121
timestamp 1683038052
transform 1 0 544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_122
timestamp 1683038052
transform 1 0 552 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1683038052
transform -1 0 656 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1683038052
transform 1 0 656 0 -1 1370
box -8 -3 104 105
use FILL  FILL_123
timestamp 1683038052
transform 1 0 752 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_24
timestamp 1683038052
transform 1 0 760 0 -1 1370
box -9 -3 26 105
use NAND2X1  NAND2X1_8
timestamp 1683038052
transform 1 0 776 0 -1 1370
box -8 -3 32 105
use FILL  FILL_128
timestamp 1683038052
transform 1 0 800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_129
timestamp 1683038052
transform 1 0 808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_130
timestamp 1683038052
transform 1 0 816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_131
timestamp 1683038052
transform 1 0 824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_132
timestamp 1683038052
transform 1 0 832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_134
timestamp 1683038052
transform 1 0 840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_136
timestamp 1683038052
transform 1 0 848 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_10
timestamp 1683038052
transform -1 0 880 0 -1 1370
box -8 -3 32 105
use FILL  FILL_137
timestamp 1683038052
transform 1 0 880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_138
timestamp 1683038052
transform 1 0 888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_139
timestamp 1683038052
transform 1 0 896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_140
timestamp 1683038052
transform 1 0 904 0 -1 1370
box -8 -3 16 105
use AND2X2  AND2X2_1
timestamp 1683038052
transform 1 0 912 0 -1 1370
box -8 -3 40 105
use FILL  FILL_152
timestamp 1683038052
transform 1 0 944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_153
timestamp 1683038052
transform 1 0 952 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_26
timestamp 1683038052
transform 1 0 960 0 -1 1370
box -9 -3 26 105
use FAX1  FAX1_6
timestamp 1683038052
transform 1 0 976 0 -1 1370
box -5 -3 126 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1683038052
transform -1 0 1192 0 -1 1370
box -8 -3 104 105
use FILL  FILL_154
timestamp 1683038052
transform 1 0 1192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_156
timestamp 1683038052
transform 1 0 1200 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_28
timestamp 1683038052
transform 1 0 1208 0 -1 1370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1683038052
transform -1 0 1320 0 -1 1370
box -8 -3 104 105
use FILL  FILL_171
timestamp 1683038052
transform 1 0 1320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_172
timestamp 1683038052
transform 1 0 1328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_173
timestamp 1683038052
transform 1 0 1336 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_4
timestamp 1683038052
transform -1 0 1384 0 -1 1370
box -8 -3 46 105
use FILL  FILL_174
timestamp 1683038052
transform 1 0 1384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_175
timestamp 1683038052
transform 1 0 1392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_176
timestamp 1683038052
transform 1 0 1400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_177
timestamp 1683038052
transform 1 0 1408 0 -1 1370
box -8 -3 16 105
use FAX1  FAX1_8
timestamp 1683038052
transform -1 0 1536 0 -1 1370
box -5 -3 126 105
use INVX2  INVX2_29
timestamp 1683038052
transform 1 0 1536 0 -1 1370
box -9 -3 26 105
use FILL  FILL_178
timestamp 1683038052
transform 1 0 1552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_179
timestamp 1683038052
transform 1 0 1560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_180
timestamp 1683038052
transform 1 0 1568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_181
timestamp 1683038052
transform 1 0 1576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_182
timestamp 1683038052
transform 1 0 1584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_183
timestamp 1683038052
transform 1 0 1592 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_14
timestamp 1683038052
transform -1 0 1632 0 -1 1370
box -8 -3 34 105
use INVX2  INVX2_30
timestamp 1683038052
transform -1 0 1648 0 -1 1370
box -9 -3 26 105
use FILL  FILL_184
timestamp 1683038052
transform 1 0 1648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_185
timestamp 1683038052
transform 1 0 1656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_186
timestamp 1683038052
transform 1 0 1664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_187
timestamp 1683038052
transform 1 0 1672 0 -1 1370
box -8 -3 16 105
use FILL  FILL_188
timestamp 1683038052
transform 1 0 1680 0 -1 1370
box -8 -3 16 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_9
timestamp 1683038052
transform 1 0 1740 0 1 1270
box -10 -3 10 3
use M2_M1  M2_M1_343
timestamp 1683038052
transform 1 0 92 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1683038052
transform 1 0 68 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1683038052
transform 1 0 76 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_311
timestamp 1683038052
transform 1 0 84 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1683038052
transform 1 0 228 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1683038052
transform 1 0 252 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_272
timestamp 1683038052
transform 1 0 284 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_344
timestamp 1683038052
transform 1 0 252 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_286
timestamp 1683038052
transform 1 0 260 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_345
timestamp 1683038052
transform 1 0 276 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_287
timestamp 1683038052
transform 1 0 284 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_356
timestamp 1683038052
transform 1 0 108 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1683038052
transform 1 0 124 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1683038052
transform 1 0 164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1683038052
transform 1 0 228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1683038052
transform 1 0 236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1683038052
transform 1 0 92 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_316
timestamp 1683038052
transform 1 0 108 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_397
timestamp 1683038052
transform 1 0 140 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_326
timestamp 1683038052
transform 1 0 204 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_273
timestamp 1683038052
transform 1 0 316 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_280
timestamp 1683038052
transform 1 0 316 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_341
timestamp 1683038052
transform 1 0 332 0 1 1235
box -2 -2 2 2
use M3_M2  M3_M2_274
timestamp 1683038052
transform 1 0 364 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_275
timestamp 1683038052
transform 1 0 380 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_276
timestamp 1683038052
transform 1 0 444 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_346
timestamp 1683038052
transform 1 0 308 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1683038052
transform 1 0 316 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1683038052
transform 1 0 340 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1683038052
transform 1 0 284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1683038052
transform 1 0 292 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1683038052
transform 1 0 252 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1683038052
transform 1 0 260 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1683038052
transform 1 0 284 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_327
timestamp 1683038052
transform 1 0 268 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1683038052
transform 1 0 348 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_363
timestamp 1683038052
transform 1 0 324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1683038052
transform 1 0 308 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_301
timestamp 1683038052
transform 1 0 340 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_364
timestamp 1683038052
transform 1 0 348 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1683038052
transform 1 0 348 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_328
timestamp 1683038052
transform 1 0 316 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_329
timestamp 1683038052
transform 1 0 348 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_349
timestamp 1683038052
transform 1 0 372 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_302
timestamp 1683038052
transform 1 0 372 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_365
timestamp 1683038052
transform 1 0 380 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1683038052
transform 1 0 420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1683038052
transform 1 0 372 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1683038052
transform 1 0 460 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1683038052
transform 1 0 484 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1683038052
transform 1 0 516 0 1 1235
box -2 -2 2 2
use M3_M2  M3_M2_289
timestamp 1683038052
transform 1 0 500 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_350
timestamp 1683038052
transform 1 0 508 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_290
timestamp 1683038052
transform 1 0 516 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_351
timestamp 1683038052
transform 1 0 532 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_291
timestamp 1683038052
transform 1 0 540 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_367
timestamp 1683038052
transform 1 0 500 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1683038052
transform 1 0 516 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_303
timestamp 1683038052
transform 1 0 532 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_369
timestamp 1683038052
transform 1 0 540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1683038052
transform 1 0 540 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1683038052
transform 1 0 564 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_292
timestamp 1683038052
transform 1 0 572 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1683038052
transform 1 0 564 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_277
timestamp 1683038052
transform 1 0 604 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_407
timestamp 1683038052
transform 1 0 596 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1683038052
transform 1 0 604 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1683038052
transform 1 0 628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1683038052
transform 1 0 628 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_293
timestamp 1683038052
transform 1 0 636 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_371
timestamp 1683038052
transform 1 0 636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1683038052
transform 1 0 644 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_294
timestamp 1683038052
transform 1 0 716 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1683038052
transform 1 0 756 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_372
timestamp 1683038052
transform 1 0 652 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1683038052
transform 1 0 660 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1683038052
transform 1 0 716 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_305
timestamp 1683038052
transform 1 0 740 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_375
timestamp 1683038052
transform 1 0 756 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_312
timestamp 1683038052
transform 1 0 660 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1683038052
transform 1 0 692 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_411
timestamp 1683038052
transform 1 0 740 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_281
timestamp 1683038052
transform 1 0 804 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1683038052
transform 1 0 804 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_376
timestamp 1683038052
transform 1 0 804 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1683038052
transform 1 0 764 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1683038052
transform 1 0 772 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_317
timestamp 1683038052
transform 1 0 756 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_377
timestamp 1683038052
transform 1 0 844 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_306
timestamp 1683038052
transform 1 0 852 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_414
timestamp 1683038052
transform 1 0 828 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_330
timestamp 1683038052
transform 1 0 804 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_415
timestamp 1683038052
transform 1 0 884 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_331
timestamp 1683038052
transform 1 0 852 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1683038052
transform 1 0 908 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1683038052
transform 1 0 916 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_432
timestamp 1683038052
transform 1 0 924 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_270
timestamp 1683038052
transform 1 0 964 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_271
timestamp 1683038052
transform 1 0 980 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_378
timestamp 1683038052
transform 1 0 980 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1683038052
transform 1 0 988 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1683038052
transform 1 0 996 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1683038052
transform 1 0 964 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_314
timestamp 1683038052
transform 1 0 972 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1683038052
transform 1 0 1028 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1683038052
transform 1 0 988 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1683038052
transform 1 0 1108 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_417
timestamp 1683038052
transform 1 0 1092 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1683038052
transform 1 0 1100 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_319
timestamp 1683038052
transform 1 0 1020 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_433
timestamp 1683038052
transform 1 0 1084 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1683038052
transform 1 0 1124 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_381
timestamp 1683038052
transform 1 0 1124 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1683038052
transform 1 0 1124 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1683038052
transform 1 0 1148 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1683038052
transform 1 0 1156 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1683038052
transform 1 0 1204 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1683038052
transform 1 0 1220 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1683038052
transform 1 0 1244 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_309
timestamp 1683038052
transform 1 0 1244 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1683038052
transform 1 0 1300 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_298
timestamp 1683038052
transform 1 0 1316 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_383
timestamp 1683038052
transform 1 0 1252 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1683038052
transform 1 0 1244 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_310
timestamp 1683038052
transform 1 0 1260 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_384
timestamp 1683038052
transform 1 0 1268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1683038052
transform 1 0 1300 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1683038052
transform 1 0 1268 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_320
timestamp 1683038052
transform 1 0 1268 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1683038052
transform 1 0 1356 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_386
timestamp 1683038052
transform 1 0 1340 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_321
timestamp 1683038052
transform 1 0 1324 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1683038052
transform 1 0 1292 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1683038052
transform 1 0 1316 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_425
timestamp 1683038052
transform 1 0 1348 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1683038052
transform 1 0 1356 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_322
timestamp 1683038052
transform 1 0 1348 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_434
timestamp 1683038052
transform 1 0 1356 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_284
timestamp 1683038052
transform 1 0 1420 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_299
timestamp 1683038052
transform 1 0 1412 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_387
timestamp 1683038052
transform 1 0 1380 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1683038052
transform 1 0 1412 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1683038052
transform 1 0 1420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1683038052
transform 1 0 1388 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_323
timestamp 1683038052
transform 1 0 1388 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1683038052
transform 1 0 1476 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_390
timestamp 1683038052
transform 1 0 1476 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1683038052
transform 1 0 1436 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_334
timestamp 1683038052
transform 1 0 1372 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1683038052
transform 1 0 1388 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1683038052
transform 1 0 1412 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_278
timestamp 1683038052
transform 1 0 1508 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_391
timestamp 1683038052
transform 1 0 1540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1683038052
transform 1 0 1588 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1683038052
transform 1 0 1628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1683038052
transform 1 0 1692 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1683038052
transform 1 0 1492 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1683038052
transform 1 0 1508 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_337
timestamp 1683038052
transform 1 0 1476 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_431
timestamp 1683038052
transform 1 0 1604 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_324
timestamp 1683038052
transform 1 0 1588 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1683038052
transform 1 0 1604 0 1 1195
box -3 -3 3 3
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_10
timestamp 1683038052
transform 1 0 48 0 1 1170
box -10 -3 10 3
use NAND2X1  NAND2X1_11
timestamp 1683038052
transform 1 0 72 0 1 1170
box -8 -3 32 105
use AND2X2  AND2X2_2
timestamp 1683038052
transform 1 0 96 0 1 1170
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1683038052
transform 1 0 128 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_338
timestamp 1683038052
transform 1 0 252 0 1 1175
box -3 -3 3 3
use OAI21X1  OAI21X1_15
timestamp 1683038052
transform 1 0 224 0 1 1170
box -8 -3 34 105
use NAND2X1  NAND2X1_12
timestamp 1683038052
transform 1 0 256 0 1 1170
box -8 -3 32 105
use OAI21X1  OAI21X1_16
timestamp 1683038052
transform 1 0 280 0 1 1170
box -8 -3 34 105
use M3_M2  M3_M2_339
timestamp 1683038052
transform 1 0 348 0 1 1175
box -3 -3 3 3
use NAND3X1  NAND3X1_10
timestamp 1683038052
transform 1 0 312 0 1 1170
box -8 -3 40 105
use OAI21X1  OAI21X1_17
timestamp 1683038052
transform 1 0 344 0 1 1170
box -8 -3 34 105
use M3_M2  M3_M2_340
timestamp 1683038052
transform 1 0 460 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_19
timestamp 1683038052
transform -1 0 472 0 1 1170
box -8 -3 104 105
use FILL  FILL_189
timestamp 1683038052
transform 1 0 472 0 1 1170
box -8 -3 16 105
use FILL  FILL_190
timestamp 1683038052
transform 1 0 480 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_31
timestamp 1683038052
transform 1 0 488 0 1 1170
box -9 -3 26 105
use NAND3X1  NAND3X1_11
timestamp 1683038052
transform 1 0 504 0 1 1170
box -8 -3 40 105
use OAI21X1  OAI21X1_18
timestamp 1683038052
transform 1 0 536 0 1 1170
box -8 -3 34 105
use FILL  FILL_191
timestamp 1683038052
transform 1 0 568 0 1 1170
box -8 -3 16 105
use FILL  FILL_192
timestamp 1683038052
transform 1 0 576 0 1 1170
box -8 -3 16 105
use FILL  FILL_193
timestamp 1683038052
transform 1 0 584 0 1 1170
box -8 -3 16 105
use FILL  FILL_194
timestamp 1683038052
transform 1 0 592 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_32
timestamp 1683038052
transform 1 0 600 0 1 1170
box -9 -3 26 105
use FILL  FILL_195
timestamp 1683038052
transform 1 0 616 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_341
timestamp 1683038052
transform 1 0 652 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_33
timestamp 1683038052
transform 1 0 624 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_34
timestamp 1683038052
transform 1 0 640 0 1 1170
box -9 -3 26 105
use M3_M2  M3_M2_342
timestamp 1683038052
transform 1 0 748 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_20
timestamp 1683038052
transform -1 0 752 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_35
timestamp 1683038052
transform -1 0 768 0 1 1170
box -9 -3 26 105
use M3_M2  M3_M2_343
timestamp 1683038052
transform 1 0 828 0 1 1175
box -3 -3 3 3
use XOR2X1  XOR2X1_1
timestamp 1683038052
transform 1 0 768 0 1 1170
box -8 -3 64 105
use M3_M2  M3_M2_344
timestamp 1683038052
transform 1 0 876 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1683038052
transform 1 0 892 0 1 1175
box -3 -3 3 3
use XNOR2X1  XNOR2X1_0
timestamp 1683038052
transform -1 0 880 0 1 1170
box -8 -3 64 105
use INVX2  INVX2_36
timestamp 1683038052
transform 1 0 880 0 1 1170
box -9 -3 26 105
use FILL  FILL_196
timestamp 1683038052
transform 1 0 896 0 1 1170
box -8 -3 16 105
use FILL  FILL_197
timestamp 1683038052
transform 1 0 904 0 1 1170
box -8 -3 16 105
use FILL  FILL_198
timestamp 1683038052
transform 1 0 912 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_346
timestamp 1683038052
transform 1 0 940 0 1 1175
box -3 -3 3 3
use OR2X1  OR2X1_0
timestamp 1683038052
transform 1 0 920 0 1 1170
box -8 -3 40 105
use FILL  FILL_199
timestamp 1683038052
transform 1 0 952 0 1 1170
box -8 -3 16 105
use FILL  FILL_200
timestamp 1683038052
transform 1 0 960 0 1 1170
box -8 -3 16 105
use FILL  FILL_201
timestamp 1683038052
transform 1 0 968 0 1 1170
box -8 -3 16 105
use FAX1  FAX1_9
timestamp 1683038052
transform 1 0 976 0 1 1170
box -5 -3 126 105
use FILL  FILL_202
timestamp 1683038052
transform 1 0 1096 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_37
timestamp 1683038052
transform 1 0 1104 0 1 1170
box -9 -3 26 105
use M3_M2  M3_M2_347
timestamp 1683038052
transform 1 0 1148 0 1 1175
box -3 -3 3 3
use OAI21X1  OAI21X1_19
timestamp 1683038052
transform -1 0 1152 0 1 1170
box -8 -3 34 105
use INVX2  INVX2_38
timestamp 1683038052
transform 1 0 1152 0 1 1170
box -9 -3 26 105
use FILL  FILL_203
timestamp 1683038052
transform 1 0 1168 0 1 1170
box -8 -3 16 105
use FILL  FILL_204
timestamp 1683038052
transform 1 0 1176 0 1 1170
box -8 -3 16 105
use FILL  FILL_205
timestamp 1683038052
transform 1 0 1184 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_348
timestamp 1683038052
transform 1 0 1204 0 1 1175
box -3 -3 3 3
use FILL  FILL_206
timestamp 1683038052
transform 1 0 1192 0 1 1170
box -8 -3 16 105
use FILL  FILL_207
timestamp 1683038052
transform 1 0 1200 0 1 1170
box -8 -3 16 105
use FILL  FILL_208
timestamp 1683038052
transform 1 0 1208 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_20
timestamp 1683038052
transform 1 0 1216 0 1 1170
box -8 -3 34 105
use INVX2  INVX2_39
timestamp 1683038052
transform -1 0 1264 0 1 1170
box -9 -3 26 105
use M3_M2  M3_M2_349
timestamp 1683038052
transform 1 0 1316 0 1 1175
box -3 -3 3 3
use XOR2X1  XOR2X1_2
timestamp 1683038052
transform 1 0 1264 0 1 1170
box -8 -3 64 105
use M3_M2  M3_M2_350
timestamp 1683038052
transform 1 0 1332 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1683038052
transform 1 0 1356 0 1 1175
box -3 -3 3 3
use AND2X2  AND2X2_3
timestamp 1683038052
transform -1 0 1352 0 1 1170
box -8 -3 40 105
use OR2X1  OR2X1_1
timestamp 1683038052
transform 1 0 1352 0 1 1170
box -8 -3 40 105
use M3_M2  M3_M2_352
timestamp 1683038052
transform 1 0 1436 0 1 1175
box -3 -3 3 3
use XOR2X1  XOR2X1_3
timestamp 1683038052
transform 1 0 1384 0 1 1170
box -8 -3 64 105
use M3_M2  M3_M2_353
timestamp 1683038052
transform 1 0 1492 0 1 1175
box -3 -3 3 3
use XNOR2X1  XNOR2X1_1
timestamp 1683038052
transform 1 0 1440 0 1 1170
box -8 -3 64 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1683038052
transform 1 0 1496 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_354
timestamp 1683038052
transform 1 0 1692 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_22
timestamp 1683038052
transform 1 0 1592 0 1 1170
box -8 -3 104 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_11
timestamp 1683038052
transform 1 0 1716 0 1 1170
box -10 -3 10 3
use M3_M2  M3_M2_355
timestamp 1683038052
transform 1 0 196 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_435
timestamp 1683038052
transform 1 0 92 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_372
timestamp 1683038052
transform 1 0 108 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1683038052
transform 1 0 140 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_436
timestamp 1683038052
transform 1 0 92 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1683038052
transform 1 0 108 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1683038052
transform 1 0 196 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1683038052
transform 1 0 68 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1683038052
transform 1 0 132 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_397
timestamp 1683038052
transform 1 0 92 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1683038052
transform 1 0 132 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1683038052
transform 1 0 140 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_439
timestamp 1683038052
transform 1 0 212 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1683038052
transform 1 0 204 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_356
timestamp 1683038052
transform 1 0 236 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_365
timestamp 1683038052
transform 1 0 308 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_357
timestamp 1683038052
transform 1 0 332 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_366
timestamp 1683038052
transform 1 0 332 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1683038052
transform 1 0 284 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1683038052
transform 1 0 324 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_440
timestamp 1683038052
transform 1 0 308 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1683038052
transform 1 0 324 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1683038052
transform 1 0 220 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1683038052
transform 1 0 228 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1683038052
transform 1 0 284 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_390
timestamp 1683038052
transform 1 0 308 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1683038052
transform 1 0 220 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1683038052
transform 1 0 356 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_442
timestamp 1683038052
transform 1 0 348 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1683038052
transform 1 0 340 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1683038052
transform 1 0 324 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_413
timestamp 1683038052
transform 1 0 252 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1683038052
transform 1 0 340 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1683038052
transform 1 0 372 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_478
timestamp 1683038052
transform 1 0 356 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_391
timestamp 1683038052
transform 1 0 364 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_359
timestamp 1683038052
transform 1 0 460 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1683038052
transform 1 0 412 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_443
timestamp 1683038052
transform 1 0 460 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1683038052
transform 1 0 412 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_392
timestamp 1683038052
transform 1 0 460 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_386
timestamp 1683038052
transform 1 0 540 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_444
timestamp 1683038052
transform 1 0 564 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_360
timestamp 1683038052
transform 1 0 604 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1683038052
transform 1 0 612 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_445
timestamp 1683038052
transform 1 0 660 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1683038052
transform 1 0 484 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1683038052
transform 1 0 540 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1683038052
transform 1 0 580 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_483
timestamp 1683038052
transform 1 0 636 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_414
timestamp 1683038052
transform 1 0 660 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_510
timestamp 1683038052
transform 1 0 676 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1683038052
transform 1 0 716 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_415
timestamp 1683038052
transform 1 0 708 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1683038052
transform 1 0 740 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_447
timestamp 1683038052
transform 1 0 740 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_410
timestamp 1683038052
transform 1 0 740 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1683038052
transform 1 0 756 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_361
timestamp 1683038052
transform 1 0 772 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_367
timestamp 1683038052
transform 1 0 820 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1683038052
transform 1 0 820 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_448
timestamp 1683038052
transform 1 0 812 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1683038052
transform 1 0 836 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1683038052
transform 1 0 844 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1683038052
transform 1 0 796 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1683038052
transform 1 0 804 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_393
timestamp 1683038052
transform 1 0 812 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_486
timestamp 1683038052
transform 1 0 828 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_487
timestamp 1683038052
transform 1 0 852 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1683038052
transform 1 0 860 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_362
timestamp 1683038052
transform 1 0 884 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_368
timestamp 1683038052
transform 1 0 884 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_451
timestamp 1683038052
transform 1 0 876 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1683038052
transform 1 0 892 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_401
timestamp 1683038052
transform 1 0 876 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1683038052
transform 1 0 1004 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1683038052
transform 1 0 916 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1683038052
transform 1 0 956 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_453
timestamp 1683038052
transform 1 0 916 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_389
timestamp 1683038052
transform 1 0 932 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_454
timestamp 1683038052
transform 1 0 1004 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1683038052
transform 1 0 924 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1683038052
transform 1 0 956 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1683038052
transform 1 0 916 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_402
timestamp 1683038052
transform 1 0 924 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1683038052
transform 1 0 940 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1683038052
transform 1 0 1004 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_455
timestamp 1683038052
transform 1 0 1036 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1683038052
transform 1 0 1052 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1683038052
transform 1 0 1060 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1683038052
transform 1 0 1028 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_394
timestamp 1683038052
transform 1 0 1036 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_492
timestamp 1683038052
transform 1 0 1044 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_403
timestamp 1683038052
transform 1 0 1028 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1683038052
transform 1 0 1052 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1683038052
transform 1 0 1180 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1683038052
transform 1 0 1108 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_458
timestamp 1683038052
transform 1 0 1108 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_381
timestamp 1683038052
transform 1 0 1204 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_459
timestamp 1683038052
transform 1 0 1204 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_382
timestamp 1683038052
transform 1 0 1300 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_460
timestamp 1683038052
transform 1 0 1300 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1683038052
transform 1 0 1316 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1683038052
transform 1 0 1324 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1683038052
transform 1 0 1084 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_494
timestamp 1683038052
transform 1 0 1092 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1683038052
transform 1 0 1132 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1683038052
transform 1 0 1188 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1683038052
transform 1 0 1252 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1683038052
transform 1 0 1284 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1683038052
transform 1 0 1292 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1683038052
transform 1 0 1308 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_395
timestamp 1683038052
transform 1 0 1316 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1683038052
transform 1 0 1388 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_463
timestamp 1683038052
transform 1 0 1380 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1683038052
transform 1 0 1388 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1683038052
transform 1 0 1332 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1683038052
transform 1 0 1364 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_405
timestamp 1683038052
transform 1 0 1316 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1683038052
transform 1 0 1332 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1683038052
transform 1 0 1364 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_503
timestamp 1683038052
transform 1 0 1412 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_363
timestamp 1683038052
transform 1 0 1428 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_465
timestamp 1683038052
transform 1 0 1444 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1683038052
transform 1 0 1452 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_504
timestamp 1683038052
transform 1 0 1436 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_396
timestamp 1683038052
transform 1 0 1444 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_505
timestamp 1683038052
transform 1 0 1476 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_371
timestamp 1683038052
transform 1 0 1532 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_467
timestamp 1683038052
transform 1 0 1532 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1683038052
transform 1 0 1620 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1683038052
transform 1 0 1516 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1683038052
transform 1 0 1556 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1683038052
transform 1 0 1620 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_408
timestamp 1683038052
transform 1 0 1516 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_409
timestamp 1683038052
transform 1 0 1556 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_512
timestamp 1683038052
transform 1 0 1620 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_417
timestamp 1683038052
transform 1 0 1540 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1683038052
transform 1 0 1572 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1683038052
transform 1 0 1644 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_469
timestamp 1683038052
transform 1 0 1644 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_470
timestamp 1683038052
transform 1 0 1692 0 1 1135
box -2 -2 2 2
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_12
timestamp 1683038052
transform 1 0 24 0 1 1070
box -10 -3 10 3
use NOR2X1  NOR2X1_2
timestamp 1683038052
transform -1 0 96 0 -1 1170
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1683038052
transform 1 0 96 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_40
timestamp 1683038052
transform 1 0 192 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_41
timestamp 1683038052
transform 1 0 208 0 -1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_24
timestamp 1683038052
transform -1 0 320 0 -1 1170
box -8 -3 104 105
use OAI21X1  OAI21X1_21
timestamp 1683038052
transform -1 0 352 0 -1 1170
box -8 -3 34 105
use FILL  FILL_209
timestamp 1683038052
transform 1 0 352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_210
timestamp 1683038052
transform 1 0 360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_211
timestamp 1683038052
transform 1 0 368 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1683038052
transform -1 0 472 0 -1 1170
box -8 -3 104 105
use FILL  FILL_212
timestamp 1683038052
transform 1 0 472 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1683038052
transform -1 0 576 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1683038052
transform -1 0 672 0 -1 1170
box -8 -3 104 105
use FILL  FILL_213
timestamp 1683038052
transform 1 0 672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_214
timestamp 1683038052
transform 1 0 680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_215
timestamp 1683038052
transform 1 0 688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_216
timestamp 1683038052
transform 1 0 696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_217
timestamp 1683038052
transform 1 0 704 0 -1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_22
timestamp 1683038052
transform -1 0 744 0 -1 1170
box -8 -3 34 105
use FILL  FILL_218
timestamp 1683038052
transform 1 0 744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_219
timestamp 1683038052
transform 1 0 752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_220
timestamp 1683038052
transform 1 0 760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_221
timestamp 1683038052
transform 1 0 768 0 -1 1170
box -8 -3 16 105
use FILL  FILL_222
timestamp 1683038052
transform 1 0 776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_223
timestamp 1683038052
transform 1 0 784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_224
timestamp 1683038052
transform 1 0 792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_225
timestamp 1683038052
transform 1 0 800 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_5
timestamp 1683038052
transform 1 0 808 0 -1 1170
box -8 -3 46 105
use INVX2  INVX2_42
timestamp 1683038052
transform 1 0 848 0 -1 1170
box -9 -3 26 105
use FILL  FILL_226
timestamp 1683038052
transform 1 0 864 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_43
timestamp 1683038052
transform 1 0 872 0 -1 1170
box -9 -3 26 105
use M3_M2  M3_M2_419
timestamp 1683038052
transform 1 0 916 0 1 1075
box -3 -3 3 3
use OAI21X1  OAI21X1_23
timestamp 1683038052
transform 1 0 888 0 -1 1170
box -8 -3 34 105
use M3_M2  M3_M2_420
timestamp 1683038052
transform 1 0 1004 0 1 1075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_28
timestamp 1683038052
transform -1 0 1016 0 -1 1170
box -8 -3 104 105
use FILL  FILL_227
timestamp 1683038052
transform 1 0 1016 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_6
timestamp 1683038052
transform 1 0 1024 0 -1 1170
box -8 -3 46 105
use FILL  FILL_228
timestamp 1683038052
transform 1 0 1064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_229
timestamp 1683038052
transform 1 0 1072 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_44
timestamp 1683038052
transform 1 0 1080 0 -1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1683038052
transform 1 0 1096 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1683038052
transform 1 0 1192 0 -1 1170
box -8 -3 104 105
use AOI22X1  AOI22X1_7
timestamp 1683038052
transform 1 0 1288 0 -1 1170
box -8 -3 46 105
use XNOR2X1  XNOR2X1_2
timestamp 1683038052
transform 1 0 1328 0 -1 1170
box -8 -3 64 105
use FILL  FILL_230
timestamp 1683038052
transform 1 0 1384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_231
timestamp 1683038052
transform 1 0 1392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_232
timestamp 1683038052
transform 1 0 1400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_233
timestamp 1683038052
transform 1 0 1408 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_8
timestamp 1683038052
transform 1 0 1416 0 -1 1170
box -8 -3 46 105
use FILL  FILL_234
timestamp 1683038052
transform 1 0 1456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_235
timestamp 1683038052
transform 1 0 1464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_236
timestamp 1683038052
transform 1 0 1472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_237
timestamp 1683038052
transform 1 0 1480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_238
timestamp 1683038052
transform 1 0 1488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_239
timestamp 1683038052
transform 1 0 1496 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_45
timestamp 1683038052
transform 1 0 1504 0 -1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1683038052
transform 1 0 1520 0 -1 1170
box -8 -3 104 105
use OAI21X1  OAI21X1_24
timestamp 1683038052
transform -1 0 1648 0 -1 1170
box -8 -3 34 105
use INVX2  INVX2_46
timestamp 1683038052
transform -1 0 1664 0 -1 1170
box -9 -3 26 105
use FILL  FILL_240
timestamp 1683038052
transform 1 0 1664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_241
timestamp 1683038052
transform 1 0 1672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_242
timestamp 1683038052
transform 1 0 1680 0 -1 1170
box -8 -3 16 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_13
timestamp 1683038052
transform 1 0 1740 0 1 1070
box -10 -3 10 3
use M2_M1  M2_M1_516
timestamp 1683038052
transform 1 0 92 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1683038052
transform 1 0 84 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_481
timestamp 1683038052
transform 1 0 92 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_492
timestamp 1683038052
transform 1 0 84 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_427
timestamp 1683038052
transform 1 0 116 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1683038052
transform 1 0 132 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_517
timestamp 1683038052
transform 1 0 116 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1683038052
transform 1 0 132 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1683038052
transform 1 0 132 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_421
timestamp 1683038052
transform 1 0 228 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1683038052
transform 1 0 164 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1683038052
transform 1 0 204 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1683038052
transform 1 0 244 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_519
timestamp 1683038052
transform 1 0 148 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_461
timestamp 1683038052
transform 1 0 164 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_520
timestamp 1683038052
transform 1 0 204 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_521
timestamp 1683038052
transform 1 0 244 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1683038052
transform 1 0 228 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1683038052
transform 1 0 292 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1683038052
transform 1 0 284 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_482
timestamp 1683038052
transform 1 0 284 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1683038052
transform 1 0 324 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1683038052
transform 1 0 356 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1683038052
transform 1 0 412 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1683038052
transform 1 0 452 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_523
timestamp 1683038052
transform 1 0 332 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1683038052
transform 1 0 348 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1683038052
transform 1 0 356 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1683038052
transform 1 0 324 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1683038052
transform 1 0 316 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_462
timestamp 1683038052
transform 1 0 364 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_526
timestamp 1683038052
transform 1 0 412 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1683038052
transform 1 0 452 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1683038052
transform 1 0 436 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_493
timestamp 1683038052
transform 1 0 348 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_463
timestamp 1683038052
transform 1 0 476 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_528
timestamp 1683038052
transform 1 0 484 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_472
timestamp 1683038052
transform 1 0 484 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_423
timestamp 1683038052
transform 1 0 532 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1683038052
transform 1 0 500 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_529
timestamp 1683038052
transform 1 0 508 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1683038052
transform 1 0 492 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_580
timestamp 1683038052
transform 1 0 500 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1683038052
transform 1 0 516 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1683038052
transform 1 0 524 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1683038052
transform 1 0 532 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_483
timestamp 1683038052
transform 1 0 508 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1683038052
transform 1 0 516 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1683038052
transform 1 0 564 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1683038052
transform 1 0 548 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_584
timestamp 1683038052
transform 1 0 548 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_424
timestamp 1683038052
transform 1 0 580 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1683038052
transform 1 0 572 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1683038052
transform 1 0 580 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_515
timestamp 1683038052
transform 1 0 572 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1683038052
transform 1 0 580 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1683038052
transform 1 0 636 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1683038052
transform 1 0 644 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_429
timestamp 1683038052
transform 1 0 820 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1683038052
transform 1 0 796 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_531
timestamp 1683038052
transform 1 0 676 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1683038052
transform 1 0 692 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1683038052
transform 1 0 732 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_473
timestamp 1683038052
transform 1 0 676 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_587
timestamp 1683038052
transform 1 0 684 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_466
timestamp 1683038052
transform 1 0 740 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_534
timestamp 1683038052
transform 1 0 788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1683038052
transform 1 0 796 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1683038052
transform 1 0 708 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_474
timestamp 1683038052
transform 1 0 748 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_589
timestamp 1683038052
transform 1 0 796 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_436
timestamp 1683038052
transform 1 0 916 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1683038052
transform 1 0 932 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1683038052
transform 1 0 908 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_536
timestamp 1683038052
transform 1 0 860 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_467
timestamp 1683038052
transform 1 0 868 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1683038052
transform 1 0 980 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1683038052
transform 1 0 972 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_537
timestamp 1683038052
transform 1 0 908 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1683038052
transform 1 0 916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1683038052
transform 1 0 932 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1683038052
transform 1 0 948 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1683038052
transform 1 0 964 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_542
timestamp 1683038052
transform 1 0 980 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1683038052
transform 1 0 1004 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1683038052
transform 1 0 820 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_475
timestamp 1683038052
transform 1 0 860 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_591
timestamp 1683038052
transform 1 0 908 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1683038052
transform 1 0 924 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1683038052
transform 1 0 948 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1683038052
transform 1 0 956 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1683038052
transform 1 0 972 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_484
timestamp 1683038052
transform 1 0 908 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1683038052
transform 1 0 940 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1683038052
transform 1 0 836 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1683038052
transform 1 0 924 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_497
timestamp 1683038052
transform 1 0 948 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_596
timestamp 1683038052
transform 1 0 996 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1683038052
transform 1 0 1020 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1683038052
transform 1 0 1028 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_439
timestamp 1683038052
transform 1 0 1068 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1683038052
transform 1 0 1108 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1683038052
transform 1 0 1044 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1683038052
transform 1 0 1036 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1683038052
transform 1 0 1180 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1683038052
transform 1 0 1164 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1683038052
transform 1 0 1108 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1683038052
transform 1 0 1156 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_544
timestamp 1683038052
transform 1 0 1044 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1683038052
transform 1 0 1052 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1683038052
transform 1 0 1092 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1683038052
transform 1 0 1148 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1683038052
transform 1 0 1156 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_549
timestamp 1683038052
transform 1 0 1172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1683038052
transform 1 0 1188 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1683038052
transform 1 0 1196 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_486
timestamp 1683038052
transform 1 0 1036 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1683038052
transform 1 0 1052 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_599
timestamp 1683038052
transform 1 0 1068 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1683038052
transform 1 0 1156 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1683038052
transform 1 0 1180 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_477
timestamp 1683038052
transform 1 0 1196 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_487
timestamp 1683038052
transform 1 0 1180 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1683038052
transform 1 0 1220 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_552
timestamp 1683038052
transform 1 0 1220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1683038052
transform 1 0 1212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1683038052
transform 1 0 1228 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_455
timestamp 1683038052
transform 1 0 1268 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_553
timestamp 1683038052
transform 1 0 1252 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_554
timestamp 1683038052
transform 1 0 1268 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1683038052
transform 1 0 1276 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1683038052
transform 1 0 1244 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1683038052
transform 1 0 1260 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_478
timestamp 1683038052
transform 1 0 1276 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_606
timestamp 1683038052
transform 1 0 1292 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_431
timestamp 1683038052
transform 1 0 1316 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_456
timestamp 1683038052
transform 1 0 1308 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_556
timestamp 1683038052
transform 1 0 1316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1683038052
transform 1 0 1332 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1683038052
transform 1 0 1308 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_469
timestamp 1683038052
transform 1 0 1340 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1683038052
transform 1 0 1460 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1683038052
transform 1 0 1372 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1683038052
transform 1 0 1356 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_558
timestamp 1683038052
transform 1 0 1356 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1683038052
transform 1 0 1340 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1683038052
transform 1 0 1348 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_488
timestamp 1683038052
transform 1 0 1348 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1683038052
transform 1 0 1324 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_559
timestamp 1683038052
transform 1 0 1372 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1683038052
transform 1 0 1380 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1683038052
transform 1 0 1436 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1683038052
transform 1 0 1460 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_489
timestamp 1683038052
transform 1 0 1460 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1683038052
transform 1 0 1380 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1683038052
transform 1 0 1476 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_562
timestamp 1683038052
transform 1 0 1476 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_490
timestamp 1683038052
transform 1 0 1484 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_563
timestamp 1683038052
transform 1 0 1492 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_432
timestamp 1683038052
transform 1 0 1532 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1683038052
transform 1 0 1516 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_513
timestamp 1683038052
transform 1 0 1620 0 1 1035
box -2 -2 2 2
use M3_M2  M3_M2_460
timestamp 1683038052
transform 1 0 1620 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_564
timestamp 1683038052
transform 1 0 1516 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1683038052
transform 1 0 1532 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1683038052
transform 1 0 1540 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1683038052
transform 1 0 1556 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_568
timestamp 1683038052
transform 1 0 1572 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1683038052
transform 1 0 1596 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_570
timestamp 1683038052
transform 1 0 1612 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1683038052
transform 1 0 1500 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_479
timestamp 1683038052
transform 1 0 1532 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_612
timestamp 1683038052
transform 1 0 1540 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1683038052
transform 1 0 1548 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1683038052
transform 1 0 1564 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_480
timestamp 1683038052
transform 1 0 1572 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_615
timestamp 1683038052
transform 1 0 1580 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1683038052
transform 1 0 1604 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1683038052
transform 1 0 1620 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1683038052
transform 1 0 1636 0 1 1035
box -2 -2 2 2
use M3_M2  M3_M2_491
timestamp 1683038052
transform 1 0 1652 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_571
timestamp 1683038052
transform 1 0 1660 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_470
timestamp 1683038052
transform 1 0 1668 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_618
timestamp 1683038052
transform 1 0 1668 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_471
timestamp 1683038052
transform 1 0 1756 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_572
timestamp 1683038052
transform 1 0 1764 0 1 1015
box -2 -2 2 2
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_14
timestamp 1683038052
transform 1 0 48 0 1 970
box -10 -3 10 3
use FILL  FILL_243
timestamp 1683038052
transform 1 0 72 0 1 970
box -8 -3 16 105
use FILL  FILL_245
timestamp 1683038052
transform 1 0 80 0 1 970
box -8 -3 16 105
use FILL  FILL_247
timestamp 1683038052
transform 1 0 88 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_9
timestamp 1683038052
transform 1 0 96 0 1 970
box -8 -3 46 105
use FILL  FILL_249
timestamp 1683038052
transform 1 0 136 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1683038052
transform -1 0 240 0 1 970
box -8 -3 104 105
use INVX2  INVX2_47
timestamp 1683038052
transform -1 0 256 0 1 970
box -9 -3 26 105
use FILL  FILL_250
timestamp 1683038052
transform 1 0 256 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_500
timestamp 1683038052
transform 1 0 276 0 1 975
box -3 -3 3 3
use FILL  FILL_263
timestamp 1683038052
transform 1 0 264 0 1 970
box -8 -3 16 105
use FILL  FILL_264
timestamp 1683038052
transform 1 0 272 0 1 970
box -8 -3 16 105
use FILL  FILL_265
timestamp 1683038052
transform 1 0 280 0 1 970
box -8 -3 16 105
use OR2X1  OR2X1_2
timestamp 1683038052
transform -1 0 320 0 1 970
box -8 -3 40 105
use AND2X2  AND2X2_4
timestamp 1683038052
transform 1 0 320 0 1 970
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1683038052
transform -1 0 448 0 1 970
box -8 -3 104 105
use INVX2  INVX2_48
timestamp 1683038052
transform -1 0 464 0 1 970
box -9 -3 26 105
use FILL  FILL_266
timestamp 1683038052
transform 1 0 464 0 1 970
box -8 -3 16 105
use FILL  FILL_274
timestamp 1683038052
transform 1 0 472 0 1 970
box -8 -3 16 105
use FILL  FILL_276
timestamp 1683038052
transform 1 0 480 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_11
timestamp 1683038052
transform 1 0 488 0 1 970
box -8 -3 46 105
use INVX2  INVX2_51
timestamp 1683038052
transform 1 0 528 0 1 970
box -9 -3 26 105
use OAI21X1  OAI21X1_26
timestamp 1683038052
transform 1 0 544 0 1 970
box -8 -3 34 105
use FILL  FILL_277
timestamp 1683038052
transform 1 0 576 0 1 970
box -8 -3 16 105
use FILL  FILL_278
timestamp 1683038052
transform 1 0 584 0 1 970
box -8 -3 16 105
use FILL  FILL_279
timestamp 1683038052
transform 1 0 592 0 1 970
box -8 -3 16 105
use FILL  FILL_280
timestamp 1683038052
transform 1 0 600 0 1 970
box -8 -3 16 105
use FILL  FILL_281
timestamp 1683038052
transform 1 0 608 0 1 970
box -8 -3 16 105
use FILL  FILL_282
timestamp 1683038052
transform 1 0 616 0 1 970
box -8 -3 16 105
use FILL  FILL_283
timestamp 1683038052
transform 1 0 624 0 1 970
box -8 -3 16 105
use FILL  FILL_284
timestamp 1683038052
transform 1 0 632 0 1 970
box -8 -3 16 105
use FILL  FILL_285
timestamp 1683038052
transform 1 0 640 0 1 970
box -8 -3 16 105
use FILL  FILL_286
timestamp 1683038052
transform 1 0 648 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_501
timestamp 1683038052
transform 1 0 684 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_12
timestamp 1683038052
transform 1 0 656 0 1 970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1683038052
transform 1 0 696 0 1 970
box -8 -3 104 105
use INVX2  INVX2_52
timestamp 1683038052
transform 1 0 792 0 1 970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1683038052
transform 1 0 808 0 1 970
box -8 -3 104 105
use M3_M2  M3_M2_502
timestamp 1683038052
transform 1 0 924 0 1 975
box -3 -3 3 3
use OAI22X1  OAI22X1_3
timestamp 1683038052
transform 1 0 904 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_13
timestamp 1683038052
transform -1 0 984 0 1 970
box -8 -3 46 105
use M3_M2  M3_M2_503
timestamp 1683038052
transform 1 0 1028 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_14
timestamp 1683038052
transform 1 0 984 0 1 970
box -8 -3 46 105
use FILL  FILL_287
timestamp 1683038052
transform 1 0 1024 0 1 970
box -8 -3 16 105
use FILL  FILL_288
timestamp 1683038052
transform 1 0 1032 0 1 970
box -8 -3 16 105
use INVX2  INVX2_53
timestamp 1683038052
transform 1 0 1040 0 1 970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1683038052
transform 1 0 1056 0 1 970
box -8 -3 104 105
use AOI22X1  AOI22X1_15
timestamp 1683038052
transform -1 0 1192 0 1 970
box -8 -3 46 105
use M3_M2  M3_M2_504
timestamp 1683038052
transform 1 0 1204 0 1 975
box -3 -3 3 3
use BUFX2  BUFX2_0
timestamp 1683038052
transform 1 0 1192 0 1 970
box -5 -3 28 105
use FILL  FILL_289
timestamp 1683038052
transform 1 0 1216 0 1 970
box -8 -3 16 105
use FILL  FILL_308
timestamp 1683038052
transform 1 0 1224 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_505
timestamp 1683038052
transform 1 0 1260 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_21
timestamp 1683038052
transform -1 0 1272 0 1 970
box -8 -3 46 105
use BUFX2  BUFX2_2
timestamp 1683038052
transform 1 0 1272 0 1 970
box -5 -3 28 105
use FILL  FILL_309
timestamp 1683038052
transform 1 0 1296 0 1 970
box -8 -3 16 105
use FILL  FILL_310
timestamp 1683038052
transform 1 0 1304 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_23
timestamp 1683038052
transform 1 0 1312 0 1 970
box -8 -3 46 105
use FILL  FILL_314
timestamp 1683038052
transform 1 0 1352 0 1 970
box -8 -3 16 105
use INVX2  INVX2_55
timestamp 1683038052
transform 1 0 1360 0 1 970
box -9 -3 26 105
use M3_M2  M3_M2_506
timestamp 1683038052
transform 1 0 1468 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_38
timestamp 1683038052
transform -1 0 1472 0 1 970
box -8 -3 104 105
use FILL  FILL_315
timestamp 1683038052
transform 1 0 1472 0 1 970
box -8 -3 16 105
use FILL  FILL_329
timestamp 1683038052
transform 1 0 1480 0 1 970
box -8 -3 16 105
use FILL  FILL_331
timestamp 1683038052
transform 1 0 1488 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_24
timestamp 1683038052
transform -1 0 1536 0 1 970
box -8 -3 46 105
use M3_M2  M3_M2_507
timestamp 1683038052
transform 1 0 1548 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_25
timestamp 1683038052
transform 1 0 1536 0 1 970
box -8 -3 46 105
use M3_M2  M3_M2_508
timestamp 1683038052
transform 1 0 1604 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_26
timestamp 1683038052
transform -1 0 1616 0 1 970
box -8 -3 46 105
use FILL  FILL_332
timestamp 1683038052
transform 1 0 1616 0 1 970
box -8 -3 16 105
use FILL  FILL_333
timestamp 1683038052
transform 1 0 1624 0 1 970
box -8 -3 16 105
use FILL  FILL_342
timestamp 1683038052
transform 1 0 1632 0 1 970
box -8 -3 16 105
use FILL  FILL_344
timestamp 1683038052
transform 1 0 1640 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_509
timestamp 1683038052
transform 1 0 1660 0 1 975
box -3 -3 3 3
use INVX2  INVX2_58
timestamp 1683038052
transform 1 0 1648 0 1 970
box -9 -3 26 105
use INVX2  INVX2_59
timestamp 1683038052
transform 1 0 1664 0 1 970
box -9 -3 26 105
use FILL  FILL_346
timestamp 1683038052
transform 1 0 1680 0 1 970
box -8 -3 16 105
use M2_M1  M2_M1_661
timestamp 1683038052
transform 1 0 68 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_565
timestamp 1683038052
transform 1 0 68 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_626
timestamp 1683038052
transform 1 0 84 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_551
timestamp 1683038052
transform 1 0 100 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_627
timestamp 1683038052
transform 1 0 132 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1683038052
transform 1 0 124 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_552
timestamp 1683038052
transform 1 0 132 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_710
timestamp 1683038052
transform 1 0 148 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1683038052
transform 1 0 156 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_576
timestamp 1683038052
transform 1 0 156 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_628
timestamp 1683038052
transform 1 0 212 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_518
timestamp 1683038052
transform 1 0 236 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_629
timestamp 1683038052
transform 1 0 236 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_543
timestamp 1683038052
transform 1 0 276 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_630
timestamp 1683038052
transform 1 0 292 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1683038052
transform 1 0 268 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1683038052
transform 1 0 276 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1683038052
transform 1 0 284 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_544
timestamp 1683038052
transform 1 0 332 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_510
timestamp 1683038052
transform 1 0 348 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_667
timestamp 1683038052
transform 1 0 332 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_553
timestamp 1683038052
transform 1 0 340 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_620
timestamp 1683038052
transform 1 0 452 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1683038052
transform 1 0 348 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1683038052
transform 1 0 356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1683038052
transform 1 0 364 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_577
timestamp 1683038052
transform 1 0 348 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1683038052
transform 1 0 412 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_671
timestamp 1683038052
transform 1 0 468 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_533
timestamp 1683038052
transform 1 0 476 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_631
timestamp 1683038052
transform 1 0 484 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1683038052
transform 1 0 492 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1683038052
transform 1 0 508 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1683038052
transform 1 0 516 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1683038052
transform 1 0 500 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_566
timestamp 1683038052
transform 1 0 484 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1683038052
transform 1 0 476 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1683038052
transform 1 0 516 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1683038052
transform 1 0 492 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_534
timestamp 1683038052
transform 1 0 532 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_673
timestamp 1683038052
transform 1 0 532 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_519
timestamp 1683038052
transform 1 0 548 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_674
timestamp 1683038052
transform 1 0 548 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_511
timestamp 1683038052
transform 1 0 644 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1683038052
transform 1 0 772 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1683038052
transform 1 0 692 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1683038052
transform 1 0 796 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_621
timestamp 1683038052
transform 1 0 676 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1683038052
transform 1 0 796 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1683038052
transform 1 0 684 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_636
timestamp 1683038052
transform 1 0 692 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1683038052
transform 1 0 588 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_555
timestamp 1683038052
transform 1 0 620 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_513
timestamp 1683038052
transform 1 0 828 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_637
timestamp 1683038052
transform 1 0 820 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1683038052
transform 1 0 836 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_514
timestamp 1683038052
transform 1 0 932 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_522
timestamp 1683038052
transform 1 0 924 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1683038052
transform 1 0 860 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_639
timestamp 1683038052
transform 1 0 860 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1683038052
transform 1 0 692 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1683038052
transform 1 0 708 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1683038052
transform 1 0 812 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1683038052
transform 1 0 828 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1683038052
transform 1 0 844 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_567
timestamp 1683038052
transform 1 0 588 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1683038052
transform 1 0 684 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1683038052
transform 1 0 708 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_587
timestamp 1683038052
transform 1 0 668 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1683038052
transform 1 0 820 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_556
timestamp 1683038052
transform 1 0 860 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_681
timestamp 1683038052
transform 1 0 900 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_557
timestamp 1683038052
transform 1 0 908 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1683038052
transform 1 0 972 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_640
timestamp 1683038052
transform 1 0 956 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1683038052
transform 1 0 972 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1683038052
transform 1 0 940 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1683038052
transform 1 0 948 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1683038052
transform 1 0 964 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_588
timestamp 1683038052
transform 1 0 884 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_558
timestamp 1683038052
transform 1 0 972 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1683038052
transform 1 0 988 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_685
timestamp 1683038052
transform 1 0 988 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_570
timestamp 1683038052
transform 1 0 980 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_545
timestamp 1683038052
transform 1 0 1004 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_686
timestamp 1683038052
transform 1 0 1004 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_516
timestamp 1683038052
transform 1 0 1020 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1683038052
transform 1 0 1020 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_623
timestamp 1683038052
transform 1 0 1020 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1683038052
transform 1 0 1020 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1683038052
transform 1 0 1028 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_559
timestamp 1683038052
transform 1 0 1020 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_644
timestamp 1683038052
transform 1 0 1044 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1683038052
transform 1 0 1036 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_571
timestamp 1683038052
transform 1 0 1020 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1683038052
transform 1 0 1036 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1683038052
transform 1 0 1028 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1683038052
transform 1 0 1044 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1683038052
transform 1 0 1068 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_688
timestamp 1683038052
transform 1 0 1060 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_560
timestamp 1683038052
transform 1 0 1084 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_525
timestamp 1683038052
transform 1 0 1132 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_645
timestamp 1683038052
transform 1 0 1116 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1683038052
transform 1 0 1132 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1683038052
transform 1 0 1100 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1683038052
transform 1 0 1108 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1683038052
transform 1 0 1124 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1683038052
transform 1 0 1148 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1683038052
transform 1 0 1148 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_583
timestamp 1683038052
transform 1 0 1148 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1683038052
transform 1 0 1148 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1683038052
transform 1 0 1156 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_526
timestamp 1683038052
transform 1 0 1172 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1683038052
transform 1 0 1188 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_647
timestamp 1683038052
transform 1 0 1188 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_527
timestamp 1683038052
transform 1 0 1204 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_625
timestamp 1683038052
transform 1 0 1204 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1683038052
transform 1 0 1180 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1683038052
transform 1 0 1196 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_561
timestamp 1683038052
transform 1 0 1204 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_573
timestamp 1683038052
transform 1 0 1196 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_648
timestamp 1683038052
transform 1 0 1220 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_591
timestamp 1683038052
transform 1 0 1212 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_528
timestamp 1683038052
transform 1 0 1244 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1683038052
transform 1 0 1244 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_649
timestamp 1683038052
transform 1 0 1244 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_562
timestamp 1683038052
transform 1 0 1236 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_546
timestamp 1683038052
transform 1 0 1252 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_695
timestamp 1683038052
transform 1 0 1244 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1683038052
transform 1 0 1252 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_584
timestamp 1683038052
transform 1 0 1252 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1683038052
transform 1 0 1276 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_650
timestamp 1683038052
transform 1 0 1292 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1683038052
transform 1 0 1300 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1683038052
transform 1 0 1284 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1683038052
transform 1 0 1300 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_574
timestamp 1683038052
transform 1 0 1284 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1683038052
transform 1 0 1300 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1683038052
transform 1 0 1284 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1683038052
transform 1 0 1316 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_699
timestamp 1683038052
transform 1 0 1348 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1683038052
transform 1 0 1356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1683038052
transform 1 0 1380 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1683038052
transform 1 0 1428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1683038052
transform 1 0 1452 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1683038052
transform 1 0 1460 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1683038052
transform 1 0 1476 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1683038052
transform 1 0 1492 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_539
timestamp 1683038052
transform 1 0 1524 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1683038052
transform 1 0 1556 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_548
timestamp 1683038052
transform 1 0 1540 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_702
timestamp 1683038052
transform 1 0 1524 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1683038052
transform 1 0 1540 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_704
timestamp 1683038052
transform 1 0 1556 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_593
timestamp 1683038052
transform 1 0 1524 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_530
timestamp 1683038052
transform 1 0 1572 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1683038052
transform 1 0 1564 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1683038052
transform 1 0 1556 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1683038052
transform 1 0 1596 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_541
timestamp 1683038052
transform 1 0 1588 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_542
timestamp 1683038052
transform 1 0 1612 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_656
timestamp 1683038052
transform 1 0 1588 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1683038052
transform 1 0 1596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1683038052
transform 1 0 1588 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_563
timestamp 1683038052
transform 1 0 1596 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_658
timestamp 1683038052
transform 1 0 1628 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1683038052
transform 1 0 1604 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_707
timestamp 1683038052
transform 1 0 1620 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_595
timestamp 1683038052
transform 1 0 1588 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_659
timestamp 1683038052
transform 1 0 1644 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_564
timestamp 1683038052
transform 1 0 1636 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1683038052
transform 1 0 1644 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_708
timestamp 1683038052
transform 1 0 1652 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_517
timestamp 1683038052
transform 1 0 1700 0 1 965
box -3 -3 3 3
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_15
timestamp 1683038052
transform 1 0 1716 0 1 970
box -10 -3 10 3
use M3_M2  M3_M2_532
timestamp 1683038052
transform 1 0 1692 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_549
timestamp 1683038052
transform 1 0 1668 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_660
timestamp 1683038052
transform 1 0 1676 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_550
timestamp 1683038052
transform 1 0 1700 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_709
timestamp 1683038052
transform 1 0 1692 0 1 925
box -2 -2 2 2
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_16
timestamp 1683038052
transform 1 0 24 0 1 870
box -10 -3 10 3
use FILL  FILL_244
timestamp 1683038052
transform 1 0 72 0 -1 970
box -8 -3 16 105
use FILL  FILL_246
timestamp 1683038052
transform 1 0 80 0 -1 970
box -8 -3 16 105
use FILL  FILL_248
timestamp 1683038052
transform 1 0 88 0 -1 970
box -8 -3 16 105
use FILL  FILL_251
timestamp 1683038052
transform 1 0 96 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_10
timestamp 1683038052
transform 1 0 104 0 -1 970
box -8 -3 46 105
use FILL  FILL_252
timestamp 1683038052
transform 1 0 144 0 -1 970
box -8 -3 16 105
use FILL  FILL_253
timestamp 1683038052
transform 1 0 152 0 -1 970
box -8 -3 16 105
use FILL  FILL_254
timestamp 1683038052
transform 1 0 160 0 -1 970
box -8 -3 16 105
use FILL  FILL_255
timestamp 1683038052
transform 1 0 168 0 -1 970
box -8 -3 16 105
use FILL  FILL_256
timestamp 1683038052
transform 1 0 176 0 -1 970
box -8 -3 16 105
use FILL  FILL_257
timestamp 1683038052
transform 1 0 184 0 -1 970
box -8 -3 16 105
use FILL  FILL_258
timestamp 1683038052
transform 1 0 192 0 -1 970
box -8 -3 16 105
use FILL  FILL_259
timestamp 1683038052
transform 1 0 200 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_25
timestamp 1683038052
transform -1 0 240 0 -1 970
box -8 -3 34 105
use FILL  FILL_260
timestamp 1683038052
transform 1 0 240 0 -1 970
box -8 -3 16 105
use FILL  FILL_261
timestamp 1683038052
transform 1 0 248 0 -1 970
box -8 -3 16 105
use FILL  FILL_262
timestamp 1683038052
transform 1 0 256 0 -1 970
box -8 -3 16 105
use FILL  FILL_267
timestamp 1683038052
transform 1 0 264 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_49
timestamp 1683038052
transform -1 0 288 0 -1 970
box -9 -3 26 105
use FILL  FILL_268
timestamp 1683038052
transform 1 0 288 0 -1 970
box -8 -3 16 105
use FILL  FILL_269
timestamp 1683038052
transform 1 0 296 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_50
timestamp 1683038052
transform -1 0 320 0 -1 970
box -9 -3 26 105
use FILL  FILL_270
timestamp 1683038052
transform 1 0 320 0 -1 970
box -8 -3 16 105
use FILL  FILL_271
timestamp 1683038052
transform 1 0 328 0 -1 970
box -8 -3 16 105
use FILL  FILL_272
timestamp 1683038052
transform 1 0 336 0 -1 970
box -8 -3 16 105
use FAX1  FAX1_10
timestamp 1683038052
transform 1 0 344 0 -1 970
box -5 -3 126 105
use FILL  FILL_273
timestamp 1683038052
transform 1 0 464 0 -1 970
box -8 -3 16 105
use FILL  FILL_275
timestamp 1683038052
transform 1 0 472 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_16
timestamp 1683038052
transform 1 0 480 0 -1 970
box -8 -3 46 105
use FILL  FILL_290
timestamp 1683038052
transform 1 0 520 0 -1 970
box -8 -3 16 105
use FILL  FILL_291
timestamp 1683038052
transform 1 0 528 0 -1 970
box -8 -3 16 105
use FILL  FILL_292
timestamp 1683038052
transform 1 0 536 0 -1 970
box -8 -3 16 105
use FILL  FILL_293
timestamp 1683038052
transform 1 0 544 0 -1 970
box -8 -3 16 105
use FILL  FILL_294
timestamp 1683038052
transform 1 0 552 0 -1 970
box -8 -3 16 105
use FILL  FILL_295
timestamp 1683038052
transform 1 0 560 0 -1 970
box -8 -3 16 105
use FAX1  FAX1_11
timestamp 1683038052
transform 1 0 568 0 -1 970
box -5 -3 126 105
use FAX1  FAX1_12
timestamp 1683038052
transform 1 0 688 0 -1 970
box -5 -3 126 105
use AOI22X1  AOI22X1_17
timestamp 1683038052
transform 1 0 808 0 -1 970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1683038052
transform 1 0 848 0 -1 970
box -8 -3 104 105
use AOI22X1  AOI22X1_18
timestamp 1683038052
transform -1 0 984 0 -1 970
box -8 -3 46 105
use FILL  FILL_296
timestamp 1683038052
transform 1 0 984 0 -1 970
box -8 -3 16 105
use FILL  FILL_297
timestamp 1683038052
transform 1 0 992 0 -1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_3
timestamp 1683038052
transform -1 0 1024 0 -1 970
box -8 -3 32 105
use INVX2  INVX2_54
timestamp 1683038052
transform 1 0 1024 0 -1 970
box -9 -3 26 105
use BUFX2  BUFX2_1
timestamp 1683038052
transform -1 0 1064 0 -1 970
box -5 -3 28 105
use FILL  FILL_298
timestamp 1683038052
transform 1 0 1064 0 -1 970
box -8 -3 16 105
use FILL  FILL_299
timestamp 1683038052
transform 1 0 1072 0 -1 970
box -8 -3 16 105
use FILL  FILL_300
timestamp 1683038052
transform 1 0 1080 0 -1 970
box -8 -3 16 105
use FILL  FILL_301
timestamp 1683038052
transform 1 0 1088 0 -1 970
box -8 -3 16 105
use FILL  FILL_302
timestamp 1683038052
transform 1 0 1096 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_19
timestamp 1683038052
transform -1 0 1144 0 -1 970
box -8 -3 46 105
use FILL  FILL_303
timestamp 1683038052
transform 1 0 1144 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_597
timestamp 1683038052
transform 1 0 1164 0 1 875
box -3 -3 3 3
use FILL  FILL_304
timestamp 1683038052
transform 1 0 1152 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_20
timestamp 1683038052
transform 1 0 1160 0 -1 970
box -8 -3 46 105
use FILL  FILL_305
timestamp 1683038052
transform 1 0 1200 0 -1 970
box -8 -3 16 105
use FILL  FILL_306
timestamp 1683038052
transform 1 0 1208 0 -1 970
box -8 -3 16 105
use FILL  FILL_307
timestamp 1683038052
transform 1 0 1216 0 -1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_4
timestamp 1683038052
transform 1 0 1224 0 -1 970
box -8 -3 32 105
use FILL  FILL_311
timestamp 1683038052
transform 1 0 1248 0 -1 970
box -8 -3 16 105
use FILL  FILL_312
timestamp 1683038052
transform 1 0 1256 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_22
timestamp 1683038052
transform 1 0 1264 0 -1 970
box -8 -3 46 105
use M3_M2  M3_M2_598
timestamp 1683038052
transform 1 0 1316 0 1 875
box -3 -3 3 3
use FILL  FILL_313
timestamp 1683038052
transform 1 0 1304 0 -1 970
box -8 -3 16 105
use FILL  FILL_316
timestamp 1683038052
transform 1 0 1312 0 -1 970
box -8 -3 16 105
use FILL  FILL_317
timestamp 1683038052
transform 1 0 1320 0 -1 970
box -8 -3 16 105
use FILL  FILL_318
timestamp 1683038052
transform 1 0 1328 0 -1 970
box -8 -3 16 105
use FILL  FILL_319
timestamp 1683038052
transform 1 0 1336 0 -1 970
box -8 -3 16 105
use FILL  FILL_320
timestamp 1683038052
transform 1 0 1344 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_56
timestamp 1683038052
transform 1 0 1352 0 -1 970
box -9 -3 26 105
use FILL  FILL_321
timestamp 1683038052
transform 1 0 1368 0 -1 970
box -8 -3 16 105
use FILL  FILL_322
timestamp 1683038052
transform 1 0 1376 0 -1 970
box -8 -3 16 105
use FILL  FILL_323
timestamp 1683038052
transform 1 0 1384 0 -1 970
box -8 -3 16 105
use FILL  FILL_324
timestamp 1683038052
transform 1 0 1392 0 -1 970
box -8 -3 16 105
use FILL  FILL_325
timestamp 1683038052
transform 1 0 1400 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_57
timestamp 1683038052
transform 1 0 1408 0 -1 970
box -9 -3 26 105
use OAI21X1  OAI21X1_27
timestamp 1683038052
transform 1 0 1424 0 -1 970
box -8 -3 34 105
use FILL  FILL_326
timestamp 1683038052
transform 1 0 1456 0 -1 970
box -8 -3 16 105
use FILL  FILL_327
timestamp 1683038052
transform 1 0 1464 0 -1 970
box -8 -3 16 105
use FILL  FILL_328
timestamp 1683038052
transform 1 0 1472 0 -1 970
box -8 -3 16 105
use FILL  FILL_330
timestamp 1683038052
transform 1 0 1480 0 -1 970
box -8 -3 16 105
use FILL  FILL_334
timestamp 1683038052
transform 1 0 1488 0 -1 970
box -8 -3 16 105
use FILL  FILL_335
timestamp 1683038052
transform 1 0 1496 0 -1 970
box -8 -3 16 105
use FILL  FILL_336
timestamp 1683038052
transform 1 0 1504 0 -1 970
box -8 -3 16 105
use FILL  FILL_337
timestamp 1683038052
transform 1 0 1512 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_599
timestamp 1683038052
transform 1 0 1548 0 1 875
box -3 -3 3 3
use AOI22X1  AOI22X1_27
timestamp 1683038052
transform -1 0 1560 0 -1 970
box -8 -3 46 105
use FILL  FILL_338
timestamp 1683038052
transform 1 0 1560 0 -1 970
box -8 -3 16 105
use FILL  FILL_339
timestamp 1683038052
transform 1 0 1568 0 -1 970
box -8 -3 16 105
use FILL  FILL_340
timestamp 1683038052
transform 1 0 1576 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_600
timestamp 1683038052
transform 1 0 1620 0 1 875
box -3 -3 3 3
use AOI22X1  AOI22X1_28
timestamp 1683038052
transform -1 0 1624 0 -1 970
box -8 -3 46 105
use M3_M2  M3_M2_601
timestamp 1683038052
transform 1 0 1636 0 1 875
box -3 -3 3 3
use FILL  FILL_341
timestamp 1683038052
transform 1 0 1624 0 -1 970
box -8 -3 16 105
use FILL  FILL_343
timestamp 1683038052
transform 1 0 1632 0 -1 970
box -8 -3 16 105
use FILL  FILL_345
timestamp 1683038052
transform 1 0 1640 0 -1 970
box -8 -3 16 105
use FILL  FILL_347
timestamp 1683038052
transform 1 0 1648 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_60
timestamp 1683038052
transform 1 0 1656 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_61
timestamp 1683038052
transform 1 0 1672 0 -1 970
box -9 -3 26 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_17
timestamp 1683038052
transform 1 0 1740 0 1 870
box -10 -3 10 3
use M3_M2  M3_M2_620
timestamp 1683038052
transform 1 0 92 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_626
timestamp 1683038052
transform 1 0 68 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_604
timestamp 1683038052
transform 1 0 196 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1683038052
transform 1 0 228 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1683038052
transform 1 0 212 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1683038052
transform 1 0 212 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_712
timestamp 1683038052
transform 1 0 212 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1683038052
transform 1 0 68 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1683038052
transform 1 0 92 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1683038052
transform 1 0 108 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1683038052
transform 1 0 172 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1683038052
transform 1 0 84 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1683038052
transform 1 0 100 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_653
timestamp 1683038052
transform 1 0 172 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_719
timestamp 1683038052
transform 1 0 228 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1683038052
transform 1 0 196 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1683038052
transform 1 0 212 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_667
timestamp 1683038052
transform 1 0 108 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1683038052
transform 1 0 276 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_720
timestamp 1683038052
transform 1 0 276 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1683038052
transform 1 0 332 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1683038052
transform 1 0 340 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_627
timestamp 1683038052
transform 1 0 348 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_723
timestamp 1683038052
transform 1 0 356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1683038052
transform 1 0 236 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1683038052
transform 1 0 252 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_654
timestamp 1683038052
transform 1 0 340 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_772
timestamp 1683038052
transform 1 0 348 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_668
timestamp 1683038052
transform 1 0 356 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1683038052
transform 1 0 380 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1683038052
transform 1 0 388 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1683038052
transform 1 0 492 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1683038052
transform 1 0 364 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_724
timestamp 1683038052
transform 1 0 372 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1683038052
transform 1 0 388 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_642
timestamp 1683038052
transform 1 0 404 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1683038052
transform 1 0 524 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_726
timestamp 1683038052
transform 1 0 412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1683038052
transform 1 0 420 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1683038052
transform 1 0 428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1683038052
transform 1 0 364 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_774
timestamp 1683038052
transform 1 0 380 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_655
timestamp 1683038052
transform 1 0 388 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_775
timestamp 1683038052
transform 1 0 396 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1683038052
transform 1 0 404 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1683038052
transform 1 0 412 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_677
timestamp 1683038052
transform 1 0 364 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1683038052
transform 1 0 540 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_729
timestamp 1683038052
transform 1 0 548 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1683038052
transform 1 0 556 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1683038052
transform 1 0 564 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_644
timestamp 1683038052
transform 1 0 580 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1683038052
transform 1 0 596 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1683038052
transform 1 0 660 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_732
timestamp 1683038052
transform 1 0 668 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1683038052
transform 1 0 524 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1683038052
transform 1 0 532 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_669
timestamp 1683038052
transform 1 0 420 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_806
timestamp 1683038052
transform 1 0 516 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_656
timestamp 1683038052
transform 1 0 540 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_780
timestamp 1683038052
transform 1 0 548 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_657
timestamp 1683038052
transform 1 0 556 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_781
timestamp 1683038052
transform 1 0 660 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1683038052
transform 1 0 668 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_670
timestamp 1683038052
transform 1 0 540 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1683038052
transform 1 0 644 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_807
timestamp 1683038052
transform 1 0 652 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_678
timestamp 1683038052
transform 1 0 524 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1683038052
transform 1 0 564 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1683038052
transform 1 0 596 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1683038052
transform 1 0 652 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_733
timestamp 1683038052
transform 1 0 684 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1683038052
transform 1 0 692 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1683038052
transform 1 0 684 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_606
timestamp 1683038052
transform 1 0 820 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1683038052
transform 1 0 844 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_608
timestamp 1683038052
transform 1 0 924 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_629
timestamp 1683038052
transform 1 0 724 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_734
timestamp 1683038052
transform 1 0 708 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1683038052
transform 1 0 724 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1683038052
transform 1 0 708 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1683038052
transform 1 0 812 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1683038052
transform 1 0 884 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_737
timestamp 1683038052
transform 1 0 916 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_647
timestamp 1683038052
transform 1 0 924 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_713
timestamp 1683038052
transform 1 0 948 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_738
timestamp 1683038052
transform 1 0 932 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1683038052
transform 1 0 836 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_658
timestamp 1683038052
transform 1 0 884 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_786
timestamp 1683038052
transform 1 0 924 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_682
timestamp 1683038052
transform 1 0 836 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1683038052
transform 1 0 940 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1683038052
transform 1 0 1044 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1683038052
transform 1 0 988 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1683038052
transform 1 0 964 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_739
timestamp 1683038052
transform 1 0 980 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1683038052
transform 1 0 988 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_741
timestamp 1683038052
transform 1 0 1044 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_787
timestamp 1683038052
transform 1 0 948 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1683038052
transform 1 0 964 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1683038052
transform 1 0 956 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_672
timestamp 1683038052
transform 1 0 964 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1683038052
transform 1 0 1068 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_789
timestamp 1683038052
transform 1 0 1068 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_683
timestamp 1683038052
transform 1 0 1068 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1683038052
transform 1 0 1116 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_618
timestamp 1683038052
transform 1 0 1124 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1683038052
transform 1 0 1140 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1683038052
transform 1 0 1092 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1683038052
transform 1 0 1108 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1683038052
transform 1 0 1132 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_742
timestamp 1683038052
transform 1 0 1092 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1683038052
transform 1 0 1108 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1683038052
transform 1 0 1124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1683038052
transform 1 0 1140 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1683038052
transform 1 0 1084 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_660
timestamp 1683038052
transform 1 0 1092 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_791
timestamp 1683038052
transform 1 0 1116 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1683038052
transform 1 0 1132 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_684
timestamp 1683038052
transform 1 0 1124 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1683038052
transform 1 0 1164 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1683038052
transform 1 0 1204 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_746
timestamp 1683038052
transform 1 0 1204 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_793
timestamp 1683038052
transform 1 0 1188 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1683038052
transform 1 0 1196 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1683038052
transform 1 0 1172 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_685
timestamp 1683038052
transform 1 0 1172 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1683038052
transform 1 0 1212 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_747
timestamp 1683038052
transform 1 0 1212 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1683038052
transform 1 0 1220 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_662
timestamp 1683038052
transform 1 0 1220 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_812
timestamp 1683038052
transform 1 0 1220 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_686
timestamp 1683038052
transform 1 0 1220 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_813
timestamp 1683038052
transform 1 0 1228 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_635
timestamp 1683038052
transform 1 0 1268 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_749
timestamp 1683038052
transform 1 0 1268 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_663
timestamp 1683038052
transform 1 0 1268 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_714
timestamp 1683038052
transform 1 0 1284 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1683038052
transform 1 0 1284 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_624
timestamp 1683038052
transform 1 0 1380 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_636
timestamp 1683038052
transform 1 0 1396 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_750
timestamp 1683038052
transform 1 0 1300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1683038052
transform 1 0 1356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1683038052
transform 1 0 1396 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1683038052
transform 1 0 1404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1683038052
transform 1 0 1316 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_673
timestamp 1683038052
transform 1 0 1316 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_814
timestamp 1683038052
transform 1 0 1404 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_687
timestamp 1683038052
transform 1 0 1404 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1683038052
transform 1 0 1428 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1683038052
transform 1 0 1436 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_754
timestamp 1683038052
transform 1 0 1428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_755
timestamp 1683038052
transform 1 0 1436 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_664
timestamp 1683038052
transform 1 0 1428 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_756
timestamp 1683038052
transform 1 0 1476 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_757
timestamp 1683038052
transform 1 0 1492 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1683038052
transform 1 0 1460 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1683038052
transform 1 0 1468 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_665
timestamp 1683038052
transform 1 0 1492 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1683038052
transform 1 0 1492 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1683038052
transform 1 0 1524 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1683038052
transform 1 0 1548 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1683038052
transform 1 0 1516 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1683038052
transform 1 0 1532 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_758
timestamp 1683038052
transform 1 0 1524 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_759
timestamp 1683038052
transform 1 0 1540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1683038052
transform 1 0 1508 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1683038052
transform 1 0 1516 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_689
timestamp 1683038052
transform 1 0 1508 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1683038052
transform 1 0 1548 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_760
timestamp 1683038052
transform 1 0 1556 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_666
timestamp 1683038052
transform 1 0 1532 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1683038052
transform 1 0 1588 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1683038052
transform 1 0 1580 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1683038052
transform 1 0 1580 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_761
timestamp 1683038052
transform 1 0 1580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1683038052
transform 1 0 1596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1683038052
transform 1 0 1580 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1683038052
transform 1 0 1588 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1683038052
transform 1 0 1604 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_674
timestamp 1683038052
transform 1 0 1580 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_675
timestamp 1683038052
transform 1 0 1596 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_763
timestamp 1683038052
transform 1 0 1628 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1683038052
transform 1 0 1620 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_690
timestamp 1683038052
transform 1 0 1628 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_619
timestamp 1683038052
transform 1 0 1756 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_764
timestamp 1683038052
transform 1 0 1668 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1683038052
transform 1 0 1676 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_651
timestamp 1683038052
transform 1 0 1692 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1683038052
transform 1 0 1756 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_805
timestamp 1683038052
transform 1 0 1692 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_676
timestamp 1683038052
transform 1 0 1692 0 1 795
box -3 -3 3 3
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_18
timestamp 1683038052
transform 1 0 48 0 1 770
box -10 -3 10 3
use AOI22X1  AOI22X1_29
timestamp 1683038052
transform 1 0 72 0 1 770
box -8 -3 46 105
use M3_M2  M3_M2_691
timestamp 1683038052
transform 1 0 180 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_39
timestamp 1683038052
transform -1 0 208 0 1 770
box -8 -3 104 105
use M3_M2  M3_M2_692
timestamp 1683038052
transform 1 0 252 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_693
timestamp 1683038052
transform 1 0 276 0 1 775
box -3 -3 3 3
use OAI21X1  OAI21X1_28
timestamp 1683038052
transform -1 0 240 0 1 770
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1683038052
transform 1 0 240 0 1 770
box -8 -3 104 105
use INVX2  INVX2_62
timestamp 1683038052
transform -1 0 352 0 1 770
box -9 -3 26 105
use INVX2  INVX2_63
timestamp 1683038052
transform -1 0 368 0 1 770
box -9 -3 26 105
use M3_M2  M3_M2_694
timestamp 1683038052
transform 1 0 380 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1683038052
transform 1 0 404 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_30
timestamp 1683038052
transform 1 0 368 0 1 770
box -8 -3 46 105
use M3_M2  M3_M2_696
timestamp 1683038052
transform 1 0 428 0 1 775
box -3 -3 3 3
use FAX1  FAX1_13
timestamp 1683038052
transform 1 0 408 0 1 770
box -5 -3 126 105
use INVX2  INVX2_64
timestamp 1683038052
transform 1 0 528 0 1 770
box -9 -3 26 105
use FAX1  FAX1_14
timestamp 1683038052
transform 1 0 544 0 1 770
box -5 -3 126 105
use NOR2X1  NOR2X1_5
timestamp 1683038052
transform -1 0 688 0 1 770
box -8 -3 32 105
use INVX2  INVX2_65
timestamp 1683038052
transform 1 0 688 0 1 770
box -9 -3 26 105
use FAX1  FAX1_15
timestamp 1683038052
transform 1 0 704 0 1 770
box -5 -3 126 105
use M3_M2  M3_M2_697
timestamp 1683038052
transform 1 0 924 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_41
timestamp 1683038052
transform 1 0 824 0 1 770
box -8 -3 104 105
use OAI21X1  OAI21X1_29
timestamp 1683038052
transform 1 0 920 0 1 770
box -8 -3 34 105
use OR2X2  OR2X2_0
timestamp 1683038052
transform 1 0 952 0 1 770
box -7 -3 35 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1683038052
transform -1 0 1080 0 1 770
box -8 -3 104 105
use FILL  FILL_348
timestamp 1683038052
transform 1 0 1080 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_31
timestamp 1683038052
transform -1 0 1128 0 1 770
box -8 -3 46 105
use M3_M2  M3_M2_698
timestamp 1683038052
transform 1 0 1156 0 1 775
box -3 -3 3 3
use NAND2X1  NAND2X1_13
timestamp 1683038052
transform 1 0 1128 0 1 770
box -8 -3 32 105
use FILL  FILL_349
timestamp 1683038052
transform 1 0 1152 0 1 770
box -8 -3 16 105
use FILL  FILL_350
timestamp 1683038052
transform 1 0 1160 0 1 770
box -8 -3 16 105
use AOI21X1  AOI21X1_3
timestamp 1683038052
transform -1 0 1200 0 1 770
box -7 -3 39 105
use M3_M2  M3_M2_699
timestamp 1683038052
transform 1 0 1220 0 1 775
box -3 -3 3 3
use INVX2  INVX2_66
timestamp 1683038052
transform 1 0 1200 0 1 770
box -9 -3 26 105
use FILL  FILL_351
timestamp 1683038052
transform 1 0 1216 0 1 770
box -8 -3 16 105
use FILL  FILL_375
timestamp 1683038052
transform 1 0 1224 0 1 770
box -8 -3 16 105
use FILL  FILL_377
timestamp 1683038052
transform 1 0 1232 0 1 770
box -8 -3 16 105
use AOI21X1  AOI21X1_4
timestamp 1683038052
transform -1 0 1272 0 1 770
box -7 -3 39 105
use FILL  FILL_378
timestamp 1683038052
transform 1 0 1272 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_700
timestamp 1683038052
transform 1 0 1292 0 1 775
box -3 -3 3 3
use FILL  FILL_379
timestamp 1683038052
transform 1 0 1280 0 1 770
box -8 -3 16 105
use INVX2  INVX2_74
timestamp 1683038052
transform 1 0 1288 0 1 770
box -9 -3 26 105
use M3_M2  M3_M2_701
timestamp 1683038052
transform 1 0 1364 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_46
timestamp 1683038052
transform 1 0 1304 0 1 770
box -8 -3 104 105
use AOI21X1  AOI21X1_5
timestamp 1683038052
transform -1 0 1432 0 1 770
box -7 -3 39 105
use FILL  FILL_380
timestamp 1683038052
transform 1 0 1432 0 1 770
box -8 -3 16 105
use FILL  FILL_381
timestamp 1683038052
transform 1 0 1440 0 1 770
box -8 -3 16 105
use FILL  FILL_382
timestamp 1683038052
transform 1 0 1448 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_702
timestamp 1683038052
transform 1 0 1468 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_33
timestamp 1683038052
transform 1 0 1456 0 1 770
box -8 -3 46 105
use FILL  FILL_383
timestamp 1683038052
transform 1 0 1496 0 1 770
box -8 -3 16 105
use FILL  FILL_384
timestamp 1683038052
transform 1 0 1504 0 1 770
box -8 -3 16 105
use FILL  FILL_385
timestamp 1683038052
transform 1 0 1512 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_34
timestamp 1683038052
transform 1 0 1520 0 1 770
box -8 -3 46 105
use FILL  FILL_386
timestamp 1683038052
transform 1 0 1560 0 1 770
box -8 -3 16 105
use FILL  FILL_387
timestamp 1683038052
transform 1 0 1568 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_703
timestamp 1683038052
transform 1 0 1604 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_35
timestamp 1683038052
transform -1 0 1616 0 1 770
box -8 -3 46 105
use FILL  FILL_388
timestamp 1683038052
transform 1 0 1616 0 1 770
box -8 -3 16 105
use FILL  FILL_389
timestamp 1683038052
transform 1 0 1624 0 1 770
box -8 -3 16 105
use FILL  FILL_390
timestamp 1683038052
transform 1 0 1632 0 1 770
box -8 -3 16 105
use FILL  FILL_399
timestamp 1683038052
transform 1 0 1640 0 1 770
box -8 -3 16 105
use FILL  FILL_401
timestamp 1683038052
transform 1 0 1648 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_704
timestamp 1683038052
transform 1 0 1668 0 1 775
box -3 -3 3 3
use INVX2  INVX2_75
timestamp 1683038052
transform 1 0 1656 0 1 770
box -9 -3 26 105
use INVX2  INVX2_76
timestamp 1683038052
transform 1 0 1672 0 1 770
box -9 -3 26 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_19
timestamp 1683038052
transform 1 0 1716 0 1 770
box -10 -3 10 3
use M3_M2  M3_M2_720
timestamp 1683038052
transform 1 0 156 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_820
timestamp 1683038052
transform 1 0 156 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1683038052
transform 1 0 68 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1683038052
transform 1 0 132 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_705
timestamp 1683038052
transform 1 0 220 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_706
timestamp 1683038052
transform 1 0 236 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_711
timestamp 1683038052
transform 1 0 228 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1683038052
transform 1 0 268 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1683038052
transform 1 0 196 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_821
timestamp 1683038052
transform 1 0 180 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1683038052
transform 1 0 212 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1683038052
transform 1 0 260 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1683038052
transform 1 0 268 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_772
timestamp 1683038052
transform 1 0 260 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_707
timestamp 1683038052
transform 1 0 332 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1683038052
transform 1 0 356 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_815
timestamp 1683038052
transform 1 0 388 0 1 745
box -2 -2 2 2
use M3_M2  M3_M2_722
timestamp 1683038052
transform 1 0 412 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_816
timestamp 1683038052
transform 1 0 428 0 1 745
box -2 -2 2 2
use M3_M2  M3_M2_723
timestamp 1683038052
transform 1 0 500 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_724
timestamp 1683038052
transform 1 0 524 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_822
timestamp 1683038052
transform 1 0 396 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_735
timestamp 1683038052
transform 1 0 404 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_823
timestamp 1683038052
transform 1 0 412 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1683038052
transform 1 0 420 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1683038052
transform 1 0 284 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1683038052
transform 1 0 292 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1683038052
transform 1 0 300 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_749
timestamp 1683038052
transform 1 0 396 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_862
timestamp 1683038052
transform 1 0 404 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_755
timestamp 1683038052
transform 1 0 292 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1683038052
transform 1 0 404 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1683038052
transform 1 0 284 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1683038052
transform 1 0 524 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_750
timestamp 1683038052
transform 1 0 500 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1683038052
transform 1 0 548 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_825
timestamp 1683038052
transform 1 0 540 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1683038052
transform 1 0 516 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1683038052
transform 1 0 524 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1683038052
transform 1 0 532 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_751
timestamp 1683038052
transform 1 0 540 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1683038052
transform 1 0 532 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_817
timestamp 1683038052
transform 1 0 556 0 1 745
box -2 -2 2 2
use M3_M2  M3_M2_737
timestamp 1683038052
transform 1 0 556 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1683038052
transform 1 0 556 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1683038052
transform 1 0 572 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_826
timestamp 1683038052
transform 1 0 572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1683038052
transform 1 0 580 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_757
timestamp 1683038052
transform 1 0 580 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_818
timestamp 1683038052
transform 1 0 604 0 1 745
box -2 -2 2 2
use M3_M2  M3_M2_738
timestamp 1683038052
transform 1 0 596 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_867
timestamp 1683038052
transform 1 0 596 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1683038052
transform 1 0 636 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_752
timestamp 1683038052
transform 1 0 636 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_828
timestamp 1683038052
transform 1 0 644 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1683038052
transform 1 0 668 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_758
timestamp 1683038052
transform 1 0 660 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1683038052
transform 1 0 676 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_739
timestamp 1683038052
transform 1 0 692 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1683038052
transform 1 0 716 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_869
timestamp 1683038052
transform 1 0 708 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1683038052
transform 1 0 716 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1683038052
transform 1 0 740 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1683038052
transform 1 0 732 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1683038052
transform 1 0 740 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_784
timestamp 1683038052
transform 1 0 740 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_830
timestamp 1683038052
transform 1 0 764 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_753
timestamp 1683038052
transform 1 0 764 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_831
timestamp 1683038052
transform 1 0 812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1683038052
transform 1 0 772 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1683038052
transform 1 0 796 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1683038052
transform 1 0 804 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_776
timestamp 1683038052
transform 1 0 772 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1683038052
transform 1 0 812 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_785
timestamp 1683038052
transform 1 0 804 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_876
timestamp 1683038052
transform 1 0 836 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1683038052
transform 1 0 860 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1683038052
transform 1 0 868 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_761
timestamp 1683038052
transform 1 0 860 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1683038052
transform 1 0 844 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1683038052
transform 1 0 868 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_879
timestamp 1683038052
transform 1 0 900 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1683038052
transform 1 0 916 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_726
timestamp 1683038052
transform 1 0 940 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_833
timestamp 1683038052
transform 1 0 932 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_727
timestamp 1683038052
transform 1 0 988 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_834
timestamp 1683038052
transform 1 0 988 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1683038052
transform 1 0 916 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1683038052
transform 1 0 924 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1683038052
transform 1 0 940 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1683038052
transform 1 0 964 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1683038052
transform 1 0 972 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1683038052
transform 1 0 980 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_762
timestamp 1683038052
transform 1 0 932 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1683038052
transform 1 0 964 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1683038052
transform 1 0 980 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_886
timestamp 1683038052
transform 1 0 1012 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1683038052
transform 1 0 1004 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_764
timestamp 1683038052
transform 1 0 1012 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_788
timestamp 1683038052
transform 1 0 1012 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_709
timestamp 1683038052
transform 1 0 1116 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_835
timestamp 1683038052
transform 1 0 1124 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1683038052
transform 1 0 1100 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_778
timestamp 1683038052
transform 1 0 1100 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1683038052
transform 1 0 1124 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1683038052
transform 1 0 1156 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_836
timestamp 1683038052
transform 1 0 1148 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1683038052
transform 1 0 1140 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_765
timestamp 1683038052
transform 1 0 1148 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1683038052
transform 1 0 1140 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1683038052
transform 1 0 1180 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_729
timestamp 1683038052
transform 1 0 1196 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_837
timestamp 1683038052
transform 1 0 1180 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_741
timestamp 1683038052
transform 1 0 1188 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_889
timestamp 1683038052
transform 1 0 1172 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1683038052
transform 1 0 1188 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_754
timestamp 1683038052
transform 1 0 1196 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_910
timestamp 1683038052
transform 1 0 1164 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_780
timestamp 1683038052
transform 1 0 1156 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1683038052
transform 1 0 1188 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1683038052
transform 1 0 1172 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1683038052
transform 1 0 1188 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1683038052
transform 1 0 1164 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1683038052
transform 1 0 1212 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_819
timestamp 1683038052
transform 1 0 1212 0 1 745
box -2 -2 2 2
use M3_M2  M3_M2_710
timestamp 1683038052
transform 1 0 1228 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1683038052
transform 1 0 1228 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_838
timestamp 1683038052
transform 1 0 1228 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1683038052
transform 1 0 1220 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_781
timestamp 1683038052
transform 1 0 1220 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1683038052
transform 1 0 1244 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_717
timestamp 1683038052
transform 1 0 1292 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_718
timestamp 1683038052
transform 1 0 1308 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1683038052
transform 1 0 1316 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_839
timestamp 1683038052
transform 1 0 1268 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1683038052
transform 1 0 1276 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_742
timestamp 1683038052
transform 1 0 1284 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_841
timestamp 1683038052
transform 1 0 1292 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_743
timestamp 1683038052
transform 1 0 1300 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_842
timestamp 1683038052
transform 1 0 1308 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1683038052
transform 1 0 1316 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1683038052
transform 1 0 1276 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1683038052
transform 1 0 1300 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_767
timestamp 1683038052
transform 1 0 1284 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1683038052
transform 1 0 1300 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1683038052
transform 1 0 1324 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_894
timestamp 1683038052
transform 1 0 1324 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_719
timestamp 1683038052
transform 1 0 1340 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_895
timestamp 1683038052
transform 1 0 1332 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_791
timestamp 1683038052
transform 1 0 1332 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1683038052
transform 1 0 1364 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_844
timestamp 1683038052
transform 1 0 1364 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1683038052
transform 1 0 1380 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_732
timestamp 1683038052
transform 1 0 1524 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_846
timestamp 1683038052
transform 1 0 1484 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_745
timestamp 1683038052
transform 1 0 1500 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_847
timestamp 1683038052
transform 1 0 1508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1683038052
transform 1 0 1524 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1683038052
transform 1 0 1356 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1683038052
transform 1 0 1372 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1683038052
transform 1 0 1388 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1683038052
transform 1 0 1404 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1683038052
transform 1 0 1436 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1683038052
transform 1 0 1500 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1683038052
transform 1 0 1516 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_768
timestamp 1683038052
transform 1 0 1356 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1683038052
transform 1 0 1380 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_911
timestamp 1683038052
transform 1 0 1396 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_782
timestamp 1683038052
transform 1 0 1388 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_783
timestamp 1683038052
transform 1 0 1436 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_792
timestamp 1683038052
transform 1 0 1404 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1683038052
transform 1 0 1540 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_903
timestamp 1683038052
transform 1 0 1540 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_770
timestamp 1683038052
transform 1 0 1540 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1683038052
transform 1 0 1580 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_849
timestamp 1683038052
transform 1 0 1556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1683038052
transform 1 0 1564 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_747
timestamp 1683038052
transform 1 0 1572 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1683038052
transform 1 0 1620 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_851
timestamp 1683038052
transform 1 0 1580 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1683038052
transform 1 0 1596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1683038052
transform 1 0 1620 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1683038052
transform 1 0 1572 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1683038052
transform 1 0 1588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1683038052
transform 1 0 1596 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1683038052
transform 1 0 1612 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1683038052
transform 1 0 1628 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_771
timestamp 1683038052
transform 1 0 1596 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1683038052
transform 1 0 1692 0 1 735
box -3 -3 3 3
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_20
timestamp 1683038052
transform 1 0 24 0 1 670
box -10 -3 10 3
use M3_M2  M3_M2_797
timestamp 1683038052
transform 1 0 68 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1683038052
transform 1 0 108 0 1 675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_43
timestamp 1683038052
transform -1 0 168 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1683038052
transform 1 0 168 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_67
timestamp 1683038052
transform -1 0 280 0 -1 770
box -9 -3 26 105
use FAX1  FAX1_16
timestamp 1683038052
transform 1 0 280 0 -1 770
box -5 -3 126 105
use INVX2  INVX2_68
timestamp 1683038052
transform -1 0 416 0 -1 770
box -9 -3 26 105
use FAX1  FAX1_17
timestamp 1683038052
transform -1 0 536 0 -1 770
box -5 -3 126 105
use FILL  FILL_352
timestamp 1683038052
transform 1 0 536 0 -1 770
box -8 -3 16 105
use FILL  FILL_353
timestamp 1683038052
transform 1 0 544 0 -1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_6
timestamp 1683038052
transform 1 0 552 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_7
timestamp 1683038052
transform -1 0 600 0 -1 770
box -8 -3 32 105
use FILL  FILL_354
timestamp 1683038052
transform 1 0 600 0 -1 770
box -8 -3 16 105
use FILL  FILL_355
timestamp 1683038052
transform 1 0 608 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_69
timestamp 1683038052
transform -1 0 632 0 -1 770
box -9 -3 26 105
use FILL  FILL_356
timestamp 1683038052
transform 1 0 632 0 -1 770
box -8 -3 16 105
use FILL  FILL_357
timestamp 1683038052
transform 1 0 640 0 -1 770
box -8 -3 16 105
use FILL  FILL_358
timestamp 1683038052
transform 1 0 648 0 -1 770
box -8 -3 16 105
use FILL  FILL_359
timestamp 1683038052
transform 1 0 656 0 -1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_8
timestamp 1683038052
transform -1 0 688 0 -1 770
box -8 -3 32 105
use FILL  FILL_360
timestamp 1683038052
transform 1 0 688 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_70
timestamp 1683038052
transform -1 0 712 0 -1 770
box -9 -3 26 105
use FILL  FILL_361
timestamp 1683038052
transform 1 0 712 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_71
timestamp 1683038052
transform -1 0 736 0 -1 770
box -9 -3 26 105
use NOR2X1  NOR2X1_9
timestamp 1683038052
transform -1 0 760 0 -1 770
box -8 -3 32 105
use MUX2X1  MUX2X1_0
timestamp 1683038052
transform -1 0 808 0 -1 770
box -5 -3 53 105
use FILL  FILL_362
timestamp 1683038052
transform 1 0 808 0 -1 770
box -8 -3 16 105
use FILL  FILL_363
timestamp 1683038052
transform 1 0 816 0 -1 770
box -8 -3 16 105
use MUX2X1  MUX2X1_1
timestamp 1683038052
transform -1 0 872 0 -1 770
box -5 -3 53 105
use FILL  FILL_364
timestamp 1683038052
transform 1 0 872 0 -1 770
box -8 -3 16 105
use FILL  FILL_365
timestamp 1683038052
transform 1 0 880 0 -1 770
box -8 -3 16 105
use FILL  FILL_366
timestamp 1683038052
transform 1 0 888 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_72
timestamp 1683038052
transform -1 0 912 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_73
timestamp 1683038052
transform 1 0 912 0 -1 770
box -9 -3 26 105
use MUX2X1  MUX2X1_2
timestamp 1683038052
transform -1 0 976 0 -1 770
box -5 -3 53 105
use FILL  FILL_367
timestamp 1683038052
transform 1 0 976 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_14
timestamp 1683038052
transform 1 0 984 0 -1 770
box -8 -3 32 105
use FILL  FILL_368
timestamp 1683038052
transform 1 0 1008 0 -1 770
box -8 -3 16 105
use FILL  FILL_369
timestamp 1683038052
transform 1 0 1016 0 -1 770
box -8 -3 16 105
use FILL  FILL_370
timestamp 1683038052
transform 1 0 1024 0 -1 770
box -8 -3 16 105
use FILL  FILL_371
timestamp 1683038052
transform 1 0 1032 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1683038052
transform -1 0 1136 0 -1 770
box -8 -3 104 105
use FILL  FILL_372
timestamp 1683038052
transform 1 0 1136 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_15
timestamp 1683038052
transform 1 0 1144 0 -1 770
box -8 -3 32 105
use AOI22X1  AOI22X1_32
timestamp 1683038052
transform -1 0 1208 0 -1 770
box -8 -3 46 105
use FILL  FILL_373
timestamp 1683038052
transform 1 0 1208 0 -1 770
box -8 -3 16 105
use FILL  FILL_374
timestamp 1683038052
transform 1 0 1216 0 -1 770
box -8 -3 16 105
use FILL  FILL_376
timestamp 1683038052
transform 1 0 1224 0 -1 770
box -8 -3 16 105
use FILL  FILL_391
timestamp 1683038052
transform 1 0 1232 0 -1 770
box -8 -3 16 105
use FILL  FILL_392
timestamp 1683038052
transform 1 0 1240 0 -1 770
box -8 -3 16 105
use FILL  FILL_393
timestamp 1683038052
transform 1 0 1248 0 -1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_10
timestamp 1683038052
transform 1 0 1256 0 -1 770
box -8 -3 32 105
use AOI22X1  AOI22X1_36
timestamp 1683038052
transform 1 0 1280 0 -1 770
box -8 -3 46 105
use FILL  FILL_394
timestamp 1683038052
transform 1 0 1320 0 -1 770
box -8 -3 16 105
use FILL  FILL_395
timestamp 1683038052
transform 1 0 1328 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_37
timestamp 1683038052
transform -1 0 1376 0 -1 770
box -8 -3 46 105
use NAND2X1  NAND2X1_16
timestamp 1683038052
transform 1 0 1376 0 -1 770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1683038052
transform -1 0 1496 0 -1 770
box -8 -3 104 105
use AOI22X1  AOI22X1_38
timestamp 1683038052
transform -1 0 1536 0 -1 770
box -8 -3 46 105
use FILL  FILL_396
timestamp 1683038052
transform 1 0 1536 0 -1 770
box -8 -3 16 105
use FILL  FILL_397
timestamp 1683038052
transform 1 0 1544 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_39
timestamp 1683038052
transform -1 0 1592 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_40
timestamp 1683038052
transform -1 0 1632 0 -1 770
box -8 -3 46 105
use FILL  FILL_398
timestamp 1683038052
transform 1 0 1632 0 -1 770
box -8 -3 16 105
use FILL  FILL_400
timestamp 1683038052
transform 1 0 1640 0 -1 770
box -8 -3 16 105
use FILL  FILL_402
timestamp 1683038052
transform 1 0 1648 0 -1 770
box -8 -3 16 105
use FILL  FILL_403
timestamp 1683038052
transform 1 0 1656 0 -1 770
box -8 -3 16 105
use FILL  FILL_404
timestamp 1683038052
transform 1 0 1664 0 -1 770
box -8 -3 16 105
use FILL  FILL_405
timestamp 1683038052
transform 1 0 1672 0 -1 770
box -8 -3 16 105
use FILL  FILL_406
timestamp 1683038052
transform 1 0 1680 0 -1 770
box -8 -3 16 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_21
timestamp 1683038052
transform 1 0 1740 0 1 670
box -10 -3 10 3
use M3_M2  M3_M2_817
timestamp 1683038052
transform 1 0 68 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_917
timestamp 1683038052
transform 1 0 68 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1683038052
transform 1 0 84 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_854
timestamp 1683038052
transform 1 0 92 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_806
timestamp 1683038052
transform 1 0 124 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1683038052
transform 1 0 108 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_918
timestamp 1683038052
transform 1 0 124 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_832
timestamp 1683038052
transform 1 0 132 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_919
timestamp 1683038052
transform 1 0 140 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1683038052
transform 1 0 148 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1683038052
transform 1 0 116 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1683038052
transform 1 0 132 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_855
timestamp 1683038052
transform 1 0 132 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_807
timestamp 1683038052
transform 1 0 196 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_912
timestamp 1683038052
transform 1 0 196 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_833
timestamp 1683038052
transform 1 0 188 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1683038052
transform 1 0 220 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1683038052
transform 1 0 324 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_921
timestamp 1683038052
transform 1 0 220 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1683038052
transform 1 0 260 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1683038052
transform 1 0 316 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1683038052
transform 1 0 324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1683038052
transform 1 0 188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1683038052
transform 1 0 196 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_841
timestamp 1683038052
transform 1 0 204 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_965
timestamp 1683038052
transform 1 0 220 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1683038052
transform 1 0 236 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_842
timestamp 1683038052
transform 1 0 260 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1683038052
transform 1 0 276 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1683038052
transform 1 0 316 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_925
timestamp 1683038052
transform 1 0 340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1683038052
transform 1 0 332 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_845
timestamp 1683038052
transform 1 0 340 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1683038052
transform 1 0 396 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1683038052
transform 1 0 516 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_834
timestamp 1683038052
transform 1 0 364 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_926
timestamp 1683038052
transform 1 0 372 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1683038052
transform 1 0 388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_928
timestamp 1683038052
transform 1 0 492 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1683038052
transform 1 0 508 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1683038052
transform 1 0 516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1683038052
transform 1 0 356 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1683038052
transform 1 0 364 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1683038052
transform 1 0 380 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_971
timestamp 1683038052
transform 1 0 396 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_856
timestamp 1683038052
transform 1 0 364 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_972
timestamp 1683038052
transform 1 0 508 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1683038052
transform 1 0 404 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_857
timestamp 1683038052
transform 1 0 428 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1683038052
transform 1 0 492 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_973
timestamp 1683038052
transform 1 0 524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1683038052
transform 1 0 540 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_865
timestamp 1683038052
transform 1 0 540 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_931
timestamp 1683038052
transform 1 0 580 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_835
timestamp 1683038052
transform 1 0 588 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_932
timestamp 1683038052
transform 1 0 596 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1683038052
transform 1 0 604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1683038052
transform 1 0 572 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_998
timestamp 1683038052
transform 1 0 580 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_866
timestamp 1683038052
transform 1 0 564 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1683038052
transform 1 0 580 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_934
timestamp 1683038052
transform 1 0 636 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_808
timestamp 1683038052
transform 1 0 692 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1683038052
transform 1 0 684 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_935
timestamp 1683038052
transform 1 0 676 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1683038052
transform 1 0 684 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1683038052
transform 1 0 692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1683038052
transform 1 0 636 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1683038052
transform 1 0 644 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_868
timestamp 1683038052
transform 1 0 628 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1683038052
transform 1 0 708 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_977
timestamp 1683038052
transform 1 0 700 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1683038052
transform 1 0 708 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1683038052
transform 1 0 716 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_869
timestamp 1683038052
transform 1 0 716 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1683038052
transform 1 0 740 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1683038052
transform 1 0 740 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_822
timestamp 1683038052
transform 1 0 764 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_938
timestamp 1683038052
transform 1 0 732 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1683038052
transform 1 0 756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1683038052
transform 1 0 764 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_870
timestamp 1683038052
transform 1 0 756 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_979
timestamp 1683038052
transform 1 0 772 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1683038052
transform 1 0 796 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_846
timestamp 1683038052
transform 1 0 796 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_823
timestamp 1683038052
transform 1 0 852 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_942
timestamp 1683038052
transform 1 0 836 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1683038052
transform 1 0 844 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1000
timestamp 1683038052
transform 1 0 876 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_824
timestamp 1683038052
transform 1 0 908 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1683038052
transform 1 0 924 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_944
timestamp 1683038052
transform 1 0 908 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1683038052
transform 1 0 932 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_803
timestamp 1683038052
transform 1 0 988 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1683038052
transform 1 0 956 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1683038052
transform 1 0 972 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1683038052
transform 1 0 996 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_946
timestamp 1683038052
transform 1 0 956 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1683038052
transform 1 0 964 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_837
timestamp 1683038052
transform 1 0 972 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_948
timestamp 1683038052
transform 1 0 988 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1683038052
transform 1 0 996 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1683038052
transform 1 0 948 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_871
timestamp 1683038052
transform 1 0 948 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1683038052
transform 1 0 1028 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1683038052
transform 1 0 1052 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1683038052
transform 1 0 1020 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1683038052
transform 1 0 1012 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_950
timestamp 1683038052
transform 1 0 1020 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_839
timestamp 1683038052
transform 1 0 1036 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_951
timestamp 1683038052
transform 1 0 1052 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_847
timestamp 1683038052
transform 1 0 1036 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_981
timestamp 1683038052
transform 1 0 1044 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1683038052
transform 1 0 1076 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_859
timestamp 1683038052
transform 1 0 1076 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_953
timestamp 1683038052
transform 1 0 1140 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_848
timestamp 1683038052
transform 1 0 1140 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_982
timestamp 1683038052
transform 1 0 1164 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1683038052
transform 1 0 1180 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_860
timestamp 1683038052
transform 1 0 1180 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1683038052
transform 1 0 1332 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_913
timestamp 1683038052
transform 1 0 1244 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_984
timestamp 1683038052
transform 1 0 1220 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_849
timestamp 1683038052
transform 1 0 1236 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1683038052
transform 1 0 1292 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1683038052
transform 1 0 1308 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_954
timestamp 1683038052
transform 1 0 1252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1683038052
transform 1 0 1308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1683038052
transform 1 0 1244 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_872
timestamp 1683038052
transform 1 0 1220 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1683038052
transform 1 0 1308 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_986
timestamp 1683038052
transform 1 0 1332 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1683038052
transform 1 0 1348 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_861
timestamp 1683038052
transform 1 0 1252 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_862
timestamp 1683038052
transform 1 0 1348 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_816
timestamp 1683038052
transform 1 0 1364 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_801
timestamp 1683038052
transform 1 0 1396 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_914
timestamp 1683038052
transform 1 0 1396 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_840
timestamp 1683038052
transform 1 0 1388 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_829
timestamp 1683038052
transform 1 0 1460 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_956
timestamp 1683038052
transform 1 0 1396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1683038052
transform 1 0 1404 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1683038052
transform 1 0 1460 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1683038052
transform 1 0 1372 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_851
timestamp 1683038052
transform 1 0 1388 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_989
timestamp 1683038052
transform 1 0 1396 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_873
timestamp 1683038052
transform 1 0 1372 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_852
timestamp 1683038052
transform 1 0 1460 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_990
timestamp 1683038052
transform 1 0 1484 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_863
timestamp 1683038052
transform 1 0 1396 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_874
timestamp 1683038052
transform 1 0 1404 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1683038052
transform 1 0 1500 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1683038052
transform 1 0 1516 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1683038052
transform 1 0 1548 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_959
timestamp 1683038052
transform 1 0 1548 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_991
timestamp 1683038052
transform 1 0 1508 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_992
timestamp 1683038052
transform 1 0 1524 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_853
timestamp 1683038052
transform 1 0 1540 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_993
timestamp 1683038052
transform 1 0 1548 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_864
timestamp 1683038052
transform 1 0 1516 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1683038052
transform 1 0 1508 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_915
timestamp 1683038052
transform 1 0 1556 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1683038052
transform 1 0 1580 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_876
timestamp 1683038052
transform 1 0 1556 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_916
timestamp 1683038052
transform 1 0 1612 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_995
timestamp 1683038052
transform 1 0 1628 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_805
timestamp 1683038052
transform 1 0 1700 0 1 645
box -3 -3 3 3
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_22
timestamp 1683038052
transform 1 0 48 0 1 570
box -10 -3 10 3
use FILL  FILL_407
timestamp 1683038052
transform 1 0 72 0 1 570
box -8 -3 16 105
use FILL  FILL_409
timestamp 1683038052
transform 1 0 80 0 1 570
box -8 -3 16 105
use FILL  FILL_411
timestamp 1683038052
transform 1 0 88 0 1 570
box -8 -3 16 105
use FILL  FILL_413
timestamp 1683038052
transform 1 0 96 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_41
timestamp 1683038052
transform 1 0 104 0 1 570
box -8 -3 46 105
use FILL  FILL_415
timestamp 1683038052
transform 1 0 144 0 1 570
box -8 -3 16 105
use FILL  FILL_417
timestamp 1683038052
transform 1 0 152 0 1 570
box -8 -3 16 105
use FILL  FILL_419
timestamp 1683038052
transform 1 0 160 0 1 570
box -8 -3 16 105
use FILL  FILL_421
timestamp 1683038052
transform 1 0 168 0 1 570
box -8 -3 16 105
use INVX2  INVX2_77
timestamp 1683038052
transform -1 0 192 0 1 570
box -9 -3 26 105
use OAI21X1  OAI21X1_30
timestamp 1683038052
transform -1 0 224 0 1 570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1683038052
transform 1 0 224 0 1 570
box -8 -3 104 105
use INVX2  INVX2_78
timestamp 1683038052
transform -1 0 336 0 1 570
box -9 -3 26 105
use FILL  FILL_422
timestamp 1683038052
transform 1 0 336 0 1 570
box -8 -3 16 105
use FILL  FILL_423
timestamp 1683038052
transform 1 0 344 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_877
timestamp 1683038052
transform 1 0 380 0 1 575
box -3 -3 3 3
use AOI22X1  AOI22X1_43
timestamp 1683038052
transform 1 0 352 0 1 570
box -8 -3 46 105
use FAX1  FAX1_18
timestamp 1683038052
transform -1 0 512 0 1 570
box -5 -3 126 105
use INVX2  INVX2_79
timestamp 1683038052
transform -1 0 528 0 1 570
box -9 -3 26 105
use FILL  FILL_424
timestamp 1683038052
transform 1 0 528 0 1 570
box -8 -3 16 105
use FILL  FILL_425
timestamp 1683038052
transform 1 0 536 0 1 570
box -8 -3 16 105
use FILL  FILL_426
timestamp 1683038052
transform 1 0 544 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_11
timestamp 1683038052
transform 1 0 552 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_12
timestamp 1683038052
transform 1 0 576 0 1 570
box -8 -3 32 105
use INVX2  INVX2_80
timestamp 1683038052
transform -1 0 616 0 1 570
box -9 -3 26 105
use FILL  FILL_427
timestamp 1683038052
transform 1 0 616 0 1 570
box -8 -3 16 105
use FILL  FILL_442
timestamp 1683038052
transform 1 0 624 0 1 570
box -8 -3 16 105
use FILL  FILL_444
timestamp 1683038052
transform 1 0 632 0 1 570
box -8 -3 16 105
use MUX2X1  MUX2X1_4
timestamp 1683038052
transform -1 0 688 0 1 570
box -5 -3 53 105
use NOR2X1  NOR2X1_14
timestamp 1683038052
transform -1 0 712 0 1 570
box -8 -3 32 105
use FILL  FILL_446
timestamp 1683038052
transform 1 0 712 0 1 570
box -8 -3 16 105
use MUX2X1  MUX2X1_5
timestamp 1683038052
transform -1 0 768 0 1 570
box -5 -3 53 105
use FILL  FILL_447
timestamp 1683038052
transform 1 0 768 0 1 570
box -8 -3 16 105
use FILL  FILL_448
timestamp 1683038052
transform 1 0 776 0 1 570
box -8 -3 16 105
use FILL  FILL_449
timestamp 1683038052
transform 1 0 784 0 1 570
box -8 -3 16 105
use FILL  FILL_450
timestamp 1683038052
transform 1 0 792 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_878
timestamp 1683038052
transform 1 0 836 0 1 575
box -3 -3 3 3
use MUX2X1  MUX2X1_6
timestamp 1683038052
transform -1 0 848 0 1 570
box -5 -3 53 105
use FILL  FILL_451
timestamp 1683038052
transform 1 0 848 0 1 570
box -8 -3 16 105
use FILL  FILL_452
timestamp 1683038052
transform 1 0 856 0 1 570
box -8 -3 16 105
use FILL  FILL_453
timestamp 1683038052
transform 1 0 864 0 1 570
box -8 -3 16 105
use FILL  FILL_454
timestamp 1683038052
transform 1 0 872 0 1 570
box -8 -3 16 105
use FILL  FILL_455
timestamp 1683038052
transform 1 0 880 0 1 570
box -8 -3 16 105
use FILL  FILL_456
timestamp 1683038052
transform 1 0 888 0 1 570
box -8 -3 16 105
use MUX2X1  MUX2X1_7
timestamp 1683038052
transform -1 0 944 0 1 570
box -5 -3 53 105
use FILL  FILL_457
timestamp 1683038052
transform 1 0 944 0 1 570
box -8 -3 16 105
use MUX2X1  MUX2X1_8
timestamp 1683038052
transform -1 0 1000 0 1 570
box -5 -3 53 105
use FILL  FILL_458
timestamp 1683038052
transform 1 0 1000 0 1 570
box -8 -3 16 105
use MUX2X1  MUX2X1_9
timestamp 1683038052
transform 1 0 1008 0 1 570
box -5 -3 53 105
use M3_M2  M3_M2_879
timestamp 1683038052
transform 1 0 1068 0 1 575
box -3 -3 3 3
use FILL  FILL_459
timestamp 1683038052
transform 1 0 1056 0 1 570
box -8 -3 16 105
use FILL  FILL_460
timestamp 1683038052
transform 1 0 1064 0 1 570
box -8 -3 16 105
use FILL  FILL_461
timestamp 1683038052
transform 1 0 1072 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_880
timestamp 1683038052
transform 1 0 1164 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_49
timestamp 1683038052
transform -1 0 1176 0 1 570
box -8 -3 104 105
use FILL  FILL_462
timestamp 1683038052
transform 1 0 1176 0 1 570
box -8 -3 16 105
use FILL  FILL_463
timestamp 1683038052
transform 1 0 1184 0 1 570
box -8 -3 16 105
use FILL  FILL_464
timestamp 1683038052
transform 1 0 1192 0 1 570
box -8 -3 16 105
use INVX2  INVX2_81
timestamp 1683038052
transform 1 0 1200 0 1 570
box -9 -3 26 105
use OAI21X1  OAI21X1_32
timestamp 1683038052
transform 1 0 1216 0 1 570
box -8 -3 34 105
use M3_M2  M3_M2_881
timestamp 1683038052
transform 1 0 1332 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_51
timestamp 1683038052
transform -1 0 1344 0 1 570
box -8 -3 104 105
use M3_M2  M3_M2_882
timestamp 1683038052
transform 1 0 1372 0 1 575
box -3 -3 3 3
use INVX2  INVX2_82
timestamp 1683038052
transform 1 0 1344 0 1 570
box -9 -3 26 105
use FILL  FILL_469
timestamp 1683038052
transform 1 0 1360 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_33
timestamp 1683038052
transform 1 0 1368 0 1 570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1683038052
transform -1 0 1496 0 1 570
box -8 -3 104 105
use FILL  FILL_470
timestamp 1683038052
transform 1 0 1496 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_883
timestamp 1683038052
transform 1 0 1524 0 1 575
box -3 -3 3 3
use INVX2  INVX2_83
timestamp 1683038052
transform 1 0 1504 0 1 570
box -9 -3 26 105
use OAI21X1  OAI21X1_34
timestamp 1683038052
transform 1 0 1520 0 1 570
box -8 -3 34 105
use FILL  FILL_471
timestamp 1683038052
transform 1 0 1552 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_884
timestamp 1683038052
transform 1 0 1580 0 1 575
box -3 -3 3 3
use INVX2  INVX2_84
timestamp 1683038052
transform 1 0 1560 0 1 570
box -9 -3 26 105
use OAI21X1  OAI21X1_35
timestamp 1683038052
transform 1 0 1576 0 1 570
box -8 -3 34 105
use FILL  FILL_472
timestamp 1683038052
transform 1 0 1608 0 1 570
box -8 -3 16 105
use FILL  FILL_473
timestamp 1683038052
transform 1 0 1616 0 1 570
box -8 -3 16 105
use FILL  FILL_474
timestamp 1683038052
transform 1 0 1624 0 1 570
box -8 -3 16 105
use FILL  FILL_475
timestamp 1683038052
transform 1 0 1632 0 1 570
box -8 -3 16 105
use FILL  FILL_476
timestamp 1683038052
transform 1 0 1640 0 1 570
box -8 -3 16 105
use FILL  FILL_477
timestamp 1683038052
transform 1 0 1648 0 1 570
box -8 -3 16 105
use FILL  FILL_478
timestamp 1683038052
transform 1 0 1656 0 1 570
box -8 -3 16 105
use FILL  FILL_479
timestamp 1683038052
transform 1 0 1664 0 1 570
box -8 -3 16 105
use FILL  FILL_480
timestamp 1683038052
transform 1 0 1672 0 1 570
box -8 -3 16 105
use FILL  FILL_481
timestamp 1683038052
transform 1 0 1680 0 1 570
box -8 -3 16 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_23
timestamp 1683038052
transform 1 0 1716 0 1 570
box -10 -3 10 3
use M2_M1  M2_M1_1029
timestamp 1683038052
transform 1 0 68 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_922
timestamp 1683038052
transform 1 0 68 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_1004
timestamp 1683038052
transform 1 0 116 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1683038052
transform 1 0 132 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1683038052
transform 1 0 124 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_917
timestamp 1683038052
transform 1 0 132 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1683038052
transform 1 0 132 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_1076
timestamp 1683038052
transform 1 0 148 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1683038052
transform 1 0 156 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1683038052
transform 1 0 204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1683038052
transform 1 0 228 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1683038052
transform 1 0 300 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1683038052
transform 1 0 300 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_885
timestamp 1683038052
transform 1 0 412 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1683038052
transform 1 0 516 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1683038052
transform 1 0 356 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1683038052
transform 1 0 420 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1683038052
transform 1 0 508 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1683038052
transform 1 0 548 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1001
timestamp 1683038052
transform 1 0 316 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1683038052
transform 1 0 436 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_898
timestamp 1683038052
transform 1 0 532 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1003
timestamp 1683038052
transform 1 0 548 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_892
timestamp 1683038052
transform 1 0 604 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_899
timestamp 1683038052
transform 1 0 596 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1009
timestamp 1683038052
transform 1 0 420 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1010
timestamp 1683038052
transform 1 0 428 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1011
timestamp 1683038052
transform 1 0 540 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_918
timestamp 1683038052
transform 1 0 380 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1033
timestamp 1683038052
transform 1 0 404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1683038052
transform 1 0 412 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_909
timestamp 1683038052
transform 1 0 548 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_910
timestamp 1683038052
transform 1 0 572 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1012
timestamp 1683038052
transform 1 0 580 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_919
timestamp 1683038052
transform 1 0 508 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1035
timestamp 1683038052
transform 1 0 524 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1683038052
transform 1 0 540 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1683038052
transform 1 0 572 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1683038052
transform 1 0 580 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_920
timestamp 1683038052
transform 1 0 596 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1683038052
transform 1 0 620 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1013
timestamp 1683038052
transform 1 0 620 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1683038052
transform 1 0 604 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1683038052
transform 1 0 612 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_923
timestamp 1683038052
transform 1 0 548 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_924
timestamp 1683038052
transform 1 0 572 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1683038052
transform 1 0 588 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1683038052
transform 1 0 364 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_935
timestamp 1683038052
transform 1 0 428 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_945
timestamp 1683038052
transform 1 0 372 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_946
timestamp 1683038052
transform 1 0 404 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1683038052
transform 1 0 428 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1683038052
transform 1 0 556 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1683038052
transform 1 0 580 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_893
timestamp 1683038052
transform 1 0 636 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1041
timestamp 1683038052
transform 1 0 636 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_901
timestamp 1683038052
transform 1 0 676 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_911
timestamp 1683038052
transform 1 0 684 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1014
timestamp 1683038052
transform 1 0 692 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_894
timestamp 1683038052
transform 1 0 748 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1683038052
transform 1 0 844 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1015
timestamp 1683038052
transform 1 0 748 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_912
timestamp 1683038052
transform 1 0 788 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1016
timestamp 1683038052
transform 1 0 796 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_913
timestamp 1683038052
transform 1 0 836 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1683038052
transform 1 0 916 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_1017
timestamp 1683038052
transform 1 0 844 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_914
timestamp 1683038052
transform 1 0 884 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1018
timestamp 1683038052
transform 1 0 900 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1683038052
transform 1 0 916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1683038052
transform 1 0 924 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1683038052
transform 1 0 676 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1043
timestamp 1683038052
transform 1 0 692 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1683038052
transform 1 0 700 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1683038052
transform 1 0 732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1683038052
transform 1 0 740 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1683038052
transform 1 0 756 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1683038052
transform 1 0 780 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1683038052
transform 1 0 788 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1683038052
transform 1 0 804 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1683038052
transform 1 0 828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1683038052
transform 1 0 836 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1683038052
transform 1 0 844 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1683038052
transform 1 0 876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1055
timestamp 1683038052
transform 1 0 884 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1683038052
transform 1 0 892 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1683038052
transform 1 0 908 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_926
timestamp 1683038052
transform 1 0 676 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1683038052
transform 1 0 732 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1683038052
transform 1 0 796 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1683038052
transform 1 0 844 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1683038052
transform 1 0 692 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1683038052
transform 1 0 740 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1683038052
transform 1 0 780 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_941
timestamp 1683038052
transform 1 0 804 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_1021
timestamp 1683038052
transform 1 0 988 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1683038052
transform 1 0 980 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_921
timestamp 1683038052
transform 1 0 988 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1683038052
transform 1 0 1060 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1022
timestamp 1683038052
transform 1 0 1068 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1683038052
transform 1 0 996 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1683038052
transform 1 0 1020 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1683038052
transform 1 0 1028 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1683038052
transform 1 0 1044 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1063
timestamp 1683038052
transform 1 0 1068 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_930
timestamp 1683038052
transform 1 0 1020 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_931
timestamp 1683038052
transform 1 0 1044 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1683038052
transform 1 0 1068 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_942
timestamp 1683038052
transform 1 0 1052 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1683038052
transform 1 0 1084 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1683038052
transform 1 0 1108 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1023
timestamp 1683038052
transform 1 0 1108 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1064
timestamp 1683038052
transform 1 0 1140 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1683038052
transform 1 0 1196 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_905
timestamp 1683038052
transform 1 0 1220 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1024
timestamp 1683038052
transform 1 0 1220 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_916
timestamp 1683038052
transform 1 0 1252 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1683038052
transform 1 0 1332 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1683038052
transform 1 0 1316 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1025
timestamp 1683038052
transform 1 0 1316 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_896
timestamp 1683038052
transform 1 0 1484 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_907
timestamp 1683038052
transform 1 0 1412 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1026
timestamp 1683038052
transform 1 0 1412 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_908
timestamp 1683038052
transform 1 0 1508 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1027
timestamp 1683038052
transform 1 0 1508 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_897
timestamp 1683038052
transform 1 0 1604 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1028
timestamp 1683038052
transform 1 0 1604 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1683038052
transform 1 0 1244 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1683038052
transform 1 0 1300 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1683038052
transform 1 0 1356 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1683038052
transform 1 0 1396 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1683038052
transform 1 0 1444 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1683038052
transform 1 0 1492 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1683038052
transform 1 0 1532 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1683038052
transform 1 0 1588 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1074
timestamp 1683038052
transform 1 0 1628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1683038052
transform 1 0 1700 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_948
timestamp 1683038052
transform 1 0 1292 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1683038052
transform 1 0 1332 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_943
timestamp 1683038052
transform 1 0 1508 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_944
timestamp 1683038052
transform 1 0 1604 0 1 505
box -3 -3 3 3
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_24
timestamp 1683038052
transform 1 0 24 0 1 470
box -10 -3 10 3
use M3_M2  M3_M2_950
timestamp 1683038052
transform 1 0 68 0 1 475
box -3 -3 3 3
use FILL  FILL_408
timestamp 1683038052
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_410
timestamp 1683038052
transform 1 0 80 0 -1 570
box -8 -3 16 105
use FILL  FILL_412
timestamp 1683038052
transform 1 0 88 0 -1 570
box -8 -3 16 105
use FILL  FILL_414
timestamp 1683038052
transform 1 0 96 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_42
timestamp 1683038052
transform 1 0 104 0 -1 570
box -8 -3 46 105
use M3_M2  M3_M2_951
timestamp 1683038052
transform 1 0 156 0 1 475
box -3 -3 3 3
use FILL  FILL_416
timestamp 1683038052
transform 1 0 144 0 -1 570
box -8 -3 16 105
use FILL  FILL_418
timestamp 1683038052
transform 1 0 152 0 -1 570
box -8 -3 16 105
use FILL  FILL_420
timestamp 1683038052
transform 1 0 160 0 -1 570
box -8 -3 16 105
use FILL  FILL_428
timestamp 1683038052
transform 1 0 168 0 -1 570
box -8 -3 16 105
use FILL  FILL_429
timestamp 1683038052
transform 1 0 176 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_952
timestamp 1683038052
transform 1 0 196 0 1 475
box -3 -3 3 3
use FILL  FILL_430
timestamp 1683038052
transform 1 0 184 0 -1 570
box -8 -3 16 105
use FILL  FILL_431
timestamp 1683038052
transform 1 0 192 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_953
timestamp 1683038052
transform 1 0 228 0 1 475
box -3 -3 3 3
use OAI21X1  OAI21X1_31
timestamp 1683038052
transform -1 0 232 0 -1 570
box -8 -3 34 105
use FILL  FILL_432
timestamp 1683038052
transform 1 0 232 0 -1 570
box -8 -3 16 105
use FILL  FILL_433
timestamp 1683038052
transform 1 0 240 0 -1 570
box -8 -3 16 105
use FILL  FILL_434
timestamp 1683038052
transform 1 0 248 0 -1 570
box -8 -3 16 105
use FILL  FILL_435
timestamp 1683038052
transform 1 0 256 0 -1 570
box -8 -3 16 105
use FILL  FILL_436
timestamp 1683038052
transform 1 0 264 0 -1 570
box -8 -3 16 105
use FILL  FILL_437
timestamp 1683038052
transform 1 0 272 0 -1 570
box -8 -3 16 105
use FILL  FILL_438
timestamp 1683038052
transform 1 0 280 0 -1 570
box -8 -3 16 105
use FILL  FILL_439
timestamp 1683038052
transform 1 0 288 0 -1 570
box -8 -3 16 105
use FILL  FILL_440
timestamp 1683038052
transform 1 0 296 0 -1 570
box -8 -3 16 105
use FAX1  FAX1_19
timestamp 1683038052
transform -1 0 424 0 -1 570
box -5 -3 126 105
use FAX1  FAX1_20
timestamp 1683038052
transform -1 0 544 0 -1 570
box -5 -3 126 105
use NOR2X1  NOR2X1_13
timestamp 1683038052
transform 1 0 544 0 -1 570
box -8 -3 32 105
use MUX2X1  MUX2X1_3
timestamp 1683038052
transform -1 0 616 0 -1 570
box -5 -3 53 105
use FILL  FILL_441
timestamp 1683038052
transform 1 0 616 0 -1 570
box -8 -3 16 105
use FILL  FILL_443
timestamp 1683038052
transform 1 0 624 0 -1 570
box -8 -3 16 105
use FILL  FILL_445
timestamp 1683038052
transform 1 0 632 0 -1 570
box -8 -3 16 105
use MUX2X1  MUX2X1_10
timestamp 1683038052
transform -1 0 688 0 -1 570
box -5 -3 53 105
use FILL  FILL_465
timestamp 1683038052
transform 1 0 688 0 -1 570
box -8 -3 16 105
use MUX2X1  MUX2X1_11
timestamp 1683038052
transform -1 0 744 0 -1 570
box -5 -3 53 105
use MUX2X1  MUX2X1_12
timestamp 1683038052
transform -1 0 792 0 -1 570
box -5 -3 53 105
use MUX2X1  MUX2X1_13
timestamp 1683038052
transform -1 0 840 0 -1 570
box -5 -3 53 105
use MUX2X1  MUX2X1_14
timestamp 1683038052
transform -1 0 888 0 -1 570
box -5 -3 53 105
use M3_M2  M3_M2_954
timestamp 1683038052
transform 1 0 916 0 1 475
box -3 -3 3 3
use AOI22X1  AOI22X1_44
timestamp 1683038052
transform 1 0 888 0 -1 570
box -8 -3 46 105
use XNOR2X1  XNOR2X1_3
timestamp 1683038052
transform -1 0 984 0 -1 570
box -8 -3 64 105
use MUX2X1  MUX2X1_15
timestamp 1683038052
transform -1 0 1032 0 -1 570
box -5 -3 53 105
use MUX2X1  MUX2X1_16
timestamp 1683038052
transform 1 0 1032 0 -1 570
box -5 -3 53 105
use FILL  FILL_466
timestamp 1683038052
transform 1 0 1080 0 -1 570
box -8 -3 16 105
use FILL  FILL_467
timestamp 1683038052
transform 1 0 1088 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_955
timestamp 1683038052
transform 1 0 1116 0 1 475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_50
timestamp 1683038052
transform 1 0 1096 0 -1 570
box -8 -3 104 105
use FILL  FILL_468
timestamp 1683038052
transform 1 0 1192 0 -1 570
box -8 -3 16 105
use FILL  FILL_482
timestamp 1683038052
transform 1 0 1200 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1683038052
transform 1 0 1208 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1683038052
transform 1 0 1304 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1683038052
transform 1 0 1400 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1683038052
transform 1 0 1496 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1683038052
transform 1 0 1592 0 -1 570
box -8 -3 104 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_25
timestamp 1683038052
transform 1 0 1740 0 1 470
box -10 -3 10 3
use M2_M1  M2_M1_1078
timestamp 1683038052
transform 1 0 68 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_956
timestamp 1683038052
transform 1 0 140 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_1079
timestamp 1683038052
transform 1 0 140 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1683038052
transform 1 0 164 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_964
timestamp 1683038052
transform 1 0 204 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1683038052
transform 1 0 252 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1080
timestamp 1683038052
transform 1 0 252 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_979
timestamp 1683038052
transform 1 0 292 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1081
timestamp 1683038052
transform 1 0 308 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1683038052
transform 1 0 316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1683038052
transform 1 0 228 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_957
timestamp 1683038052
transform 1 0 324 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_1083
timestamp 1683038052
transform 1 0 324 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1683038052
transform 1 0 324 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_989
timestamp 1683038052
transform 1 0 324 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1683038052
transform 1 0 316 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_1084
timestamp 1683038052
transform 1 0 364 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_980
timestamp 1683038052
transform 1 0 372 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1085
timestamp 1683038052
transform 1 0 380 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1683038052
transform 1 0 364 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1127
timestamp 1683038052
transform 1 0 372 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1683038052
transform 1 0 388 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1683038052
transform 1 0 404 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_990
timestamp 1683038052
transform 1 0 404 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1129
timestamp 1683038052
transform 1 0 420 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_966
timestamp 1683038052
transform 1 0 436 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_967
timestamp 1683038052
transform 1 0 524 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1130
timestamp 1683038052
transform 1 0 540 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_1005
timestamp 1683038052
transform 1 0 532 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1683038052
transform 1 0 556 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_1087
timestamp 1683038052
transform 1 0 556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1683038052
transform 1 0 564 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1683038052
transform 1 0 588 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1683038052
transform 1 0 548 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_959
timestamp 1683038052
transform 1 0 612 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_1090
timestamp 1683038052
transform 1 0 604 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_1006
timestamp 1683038052
transform 1 0 596 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_960
timestamp 1683038052
transform 1 0 660 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_968
timestamp 1683038052
transform 1 0 652 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_961
timestamp 1683038052
transform 1 0 732 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1683038052
transform 1 0 716 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1077
timestamp 1683038052
transform 1 0 732 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1683038052
transform 1 0 652 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1683038052
transform 1 0 660 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1683038052
transform 1 0 668 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1683038052
transform 1 0 676 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1683038052
transform 1 0 620 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1132
timestamp 1683038052
transform 1 0 628 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_991
timestamp 1683038052
transform 1 0 620 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1683038052
transform 1 0 612 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1683038052
transform 1 0 668 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_1133
timestamp 1683038052
transform 1 0 708 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1683038052
transform 1 0 716 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_992
timestamp 1683038052
transform 1 0 668 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1683038052
transform 1 0 756 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1095
timestamp 1683038052
transform 1 0 756 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1683038052
transform 1 0 764 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_986
timestamp 1683038052
transform 1 0 756 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1683038052
transform 1 0 788 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1135
timestamp 1683038052
transform 1 0 796 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1683038052
transform 1 0 812 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_1008
timestamp 1683038052
transform 1 0 812 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_962
timestamp 1683038052
transform 1 0 900 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_1097
timestamp 1683038052
transform 1 0 884 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1683038052
transform 1 0 900 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1099
timestamp 1683038052
transform 1 0 908 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1683038052
transform 1 0 924 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1683038052
transform 1 0 852 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_993
timestamp 1683038052
transform 1 0 852 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1009
timestamp 1683038052
transform 1 0 852 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1683038052
transform 1 0 924 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_1137
timestamp 1683038052
transform 1 0 932 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_994
timestamp 1683038052
transform 1 0 932 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1683038052
transform 1 0 956 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_1153
timestamp 1683038052
transform 1 0 956 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1683038052
transform 1 0 980 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_972
timestamp 1683038052
transform 1 0 1028 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1683038052
transform 1 0 1076 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_1102
timestamp 1683038052
transform 1 0 1020 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1103
timestamp 1683038052
transform 1 0 1028 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1683038052
transform 1 0 1036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1683038052
transform 1 0 1060 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1683038052
transform 1 0 1068 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_995
timestamp 1683038052
transform 1 0 1020 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1010
timestamp 1683038052
transform 1 0 1004 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_1138
timestamp 1683038052
transform 1 0 1060 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_996
timestamp 1683038052
transform 1 0 1052 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1139
timestamp 1683038052
transform 1 0 1076 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_1011
timestamp 1683038052
transform 1 0 1068 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1683038052
transform 1 0 1092 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1107
timestamp 1683038052
transform 1 0 1108 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_981
timestamp 1683038052
transform 1 0 1116 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1683038052
transform 1 0 1148 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1108
timestamp 1683038052
transform 1 0 1132 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1683038052
transform 1 0 1140 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1683038052
transform 1 0 1148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1683038052
transform 1 0 1100 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1683038052
transform 1 0 1116 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1683038052
transform 1 0 1124 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_997
timestamp 1683038052
transform 1 0 1100 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1111
timestamp 1683038052
transform 1 0 1172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1683038052
transform 1 0 1164 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_998
timestamp 1683038052
transform 1 0 1164 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1683038052
transform 1 0 1188 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1683038052
transform 1 0 1228 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_984
timestamp 1683038052
transform 1 0 1244 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1112
timestamp 1683038052
transform 1 0 1268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1683038052
transform 1 0 1220 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_999
timestamp 1683038052
transform 1 0 1212 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1145
timestamp 1683038052
transform 1 0 1244 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_1000
timestamp 1683038052
transform 1 0 1244 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1113
timestamp 1683038052
transform 1 0 1332 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1683038052
transform 1 0 1340 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1683038052
transform 1 0 1356 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_1001
timestamp 1683038052
transform 1 0 1404 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1154
timestamp 1683038052
transform 1 0 1412 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1683038052
transform 1 0 1444 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_975
timestamp 1683038052
transform 1 0 1508 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_976
timestamp 1683038052
transform 1 0 1540 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1116
timestamp 1683038052
transform 1 0 1516 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1683038052
transform 1 0 1524 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1683038052
transform 1 0 1540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1683038052
transform 1 0 1508 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1683038052
transform 1 0 1532 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1683038052
transform 1 0 1548 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_1002
timestamp 1683038052
transform 1 0 1508 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1683038052
transform 1 0 1532 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1119
timestamp 1683038052
transform 1 0 1572 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1683038052
transform 1 0 1572 0 1 385
box -2 -2 2 2
use M3_M2  M3_M2_977
timestamp 1683038052
transform 1 0 1588 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_978
timestamp 1683038052
transform 1 0 1628 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1120
timestamp 1683038052
transform 1 0 1588 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1683038052
transform 1 0 1628 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1122
timestamp 1683038052
transform 1 0 1692 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1683038052
transform 1 0 1604 0 1 405
box -2 -2 2 2
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_26
timestamp 1683038052
transform 1 0 48 0 1 370
box -10 -3 10 3
use FILL  FILL_483
timestamp 1683038052
transform 1 0 72 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1683038052
transform -1 0 176 0 1 370
box -8 -3 104 105
use FILL  FILL_484
timestamp 1683038052
transform 1 0 176 0 1 370
box -8 -3 16 105
use FILL  FILL_485
timestamp 1683038052
transform 1 0 184 0 1 370
box -8 -3 16 105
use FILL  FILL_486
timestamp 1683038052
transform 1 0 192 0 1 370
box -8 -3 16 105
use FILL  FILL_487
timestamp 1683038052
transform 1 0 200 0 1 370
box -8 -3 16 105
use FILL  FILL_488
timestamp 1683038052
transform 1 0 208 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_59
timestamp 1683038052
transform 1 0 216 0 1 370
box -8 -3 104 105
use INVX2  INVX2_85
timestamp 1683038052
transform -1 0 328 0 1 370
box -9 -3 26 105
use INVX2  INVX2_86
timestamp 1683038052
transform -1 0 344 0 1 370
box -9 -3 26 105
use FILL  FILL_489
timestamp 1683038052
transform 1 0 344 0 1 370
box -8 -3 16 105
use FILL  FILL_490
timestamp 1683038052
transform 1 0 352 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_45
timestamp 1683038052
transform -1 0 400 0 1 370
box -8 -3 46 105
use FILL  FILL_491
timestamp 1683038052
transform 1 0 400 0 1 370
box -8 -3 16 105
use FILL  FILL_492
timestamp 1683038052
transform 1 0 408 0 1 370
box -8 -3 16 105
use FILL  FILL_493
timestamp 1683038052
transform 1 0 416 0 1 370
box -8 -3 16 105
use FILL  FILL_494
timestamp 1683038052
transform 1 0 424 0 1 370
box -8 -3 16 105
use FILL  FILL_495
timestamp 1683038052
transform 1 0 432 0 1 370
box -8 -3 16 105
use FILL  FILL_496
timestamp 1683038052
transform 1 0 440 0 1 370
box -8 -3 16 105
use FILL  FILL_497
timestamp 1683038052
transform 1 0 448 0 1 370
box -8 -3 16 105
use FILL  FILL_498
timestamp 1683038052
transform 1 0 456 0 1 370
box -8 -3 16 105
use FILL  FILL_499
timestamp 1683038052
transform 1 0 464 0 1 370
box -8 -3 16 105
use INVX2  INVX2_87
timestamp 1683038052
transform -1 0 488 0 1 370
box -9 -3 26 105
use FILL  FILL_500
timestamp 1683038052
transform 1 0 488 0 1 370
box -8 -3 16 105
use FILL  FILL_501
timestamp 1683038052
transform 1 0 496 0 1 370
box -8 -3 16 105
use FILL  FILL_502
timestamp 1683038052
transform 1 0 504 0 1 370
box -8 -3 16 105
use FILL  FILL_503
timestamp 1683038052
transform 1 0 512 0 1 370
box -8 -3 16 105
use FILL  FILL_504
timestamp 1683038052
transform 1 0 520 0 1 370
box -8 -3 16 105
use FILL  FILL_505
timestamp 1683038052
transform 1 0 528 0 1 370
box -8 -3 16 105
use FILL  FILL_506
timestamp 1683038052
transform 1 0 536 0 1 370
box -8 -3 16 105
use FILL  FILL_507
timestamp 1683038052
transform 1 0 544 0 1 370
box -8 -3 16 105
use MUX2X1  MUX2X1_17
timestamp 1683038052
transform 1 0 552 0 1 370
box -5 -3 53 105
use FILL  FILL_510
timestamp 1683038052
transform 1 0 600 0 1 370
box -8 -3 16 105
use FILL  FILL_511
timestamp 1683038052
transform 1 0 608 0 1 370
box -8 -3 16 105
use MUX2X1  MUX2X1_19
timestamp 1683038052
transform -1 0 664 0 1 370
box -5 -3 53 105
use MUX2X1  MUX2X1_20
timestamp 1683038052
transform 1 0 664 0 1 370
box -5 -3 53 105
use NAND2X1  NAND2X1_17
timestamp 1683038052
transform 1 0 712 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_15
timestamp 1683038052
transform 1 0 736 0 1 370
box -8 -3 32 105
use FILL  FILL_512
timestamp 1683038052
transform 1 0 760 0 1 370
box -8 -3 16 105
use FILL  FILL_513
timestamp 1683038052
transform 1 0 768 0 1 370
box -8 -3 16 105
use FILL  FILL_514
timestamp 1683038052
transform 1 0 776 0 1 370
box -8 -3 16 105
use FILL  FILL_515
timestamp 1683038052
transform 1 0 784 0 1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_16
timestamp 1683038052
transform -1 0 816 0 1 370
box -8 -3 32 105
use FILL  FILL_516
timestamp 1683038052
transform 1 0 816 0 1 370
box -8 -3 16 105
use FILL  FILL_524
timestamp 1683038052
transform 1 0 824 0 1 370
box -8 -3 16 105
use FILL  FILL_525
timestamp 1683038052
transform 1 0 832 0 1 370
box -8 -3 16 105
use FILL  FILL_526
timestamp 1683038052
transform 1 0 840 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_1012
timestamp 1683038052
transform 1 0 892 0 1 375
box -3 -3 3 3
use XOR2X1  XOR2X1_4
timestamp 1683038052
transform 1 0 848 0 1 370
box -8 -3 64 105
use AND2X2  AND2X2_5
timestamp 1683038052
transform -1 0 936 0 1 370
box -8 -3 40 105
use INVX2  INVX2_89
timestamp 1683038052
transform 1 0 936 0 1 370
box -9 -3 26 105
use FILL  FILL_527
timestamp 1683038052
transform 1 0 952 0 1 370
box -8 -3 16 105
use FILL  FILL_528
timestamp 1683038052
transform 1 0 960 0 1 370
box -8 -3 16 105
use FILL  FILL_529
timestamp 1683038052
transform 1 0 968 0 1 370
box -8 -3 16 105
use FILL  FILL_530
timestamp 1683038052
transform 1 0 976 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_1013
timestamp 1683038052
transform 1 0 1012 0 1 375
box -3 -3 3 3
use OR2X1  OR2X1_3
timestamp 1683038052
transform 1 0 984 0 1 370
box -8 -3 40 105
use FILL  FILL_531
timestamp 1683038052
transform 1 0 1016 0 1 370
box -8 -3 16 105
use MUX2X1  MUX2X1_24
timestamp 1683038052
transform 1 0 1024 0 1 370
box -5 -3 53 105
use FILL  FILL_532
timestamp 1683038052
transform 1 0 1072 0 1 370
box -8 -3 16 105
use FILL  FILL_533
timestamp 1683038052
transform 1 0 1080 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_48
timestamp 1683038052
transform 1 0 1088 0 1 370
box -8 -3 46 105
use INVX2  INVX2_90
timestamp 1683038052
transform 1 0 1128 0 1 370
box -9 -3 26 105
use BUFX2  BUFX2_3
timestamp 1683038052
transform 1 0 1144 0 1 370
box -5 -3 28 105
use FILL  FILL_534
timestamp 1683038052
transform 1 0 1168 0 1 370
box -8 -3 16 105
use FILL  FILL_535
timestamp 1683038052
transform 1 0 1176 0 1 370
box -8 -3 16 105
use FILL  FILL_536
timestamp 1683038052
transform 1 0 1184 0 1 370
box -8 -3 16 105
use FILL  FILL_537
timestamp 1683038052
transform 1 0 1192 0 1 370
box -8 -3 16 105
use BUFX2  BUFX2_4
timestamp 1683038052
transform 1 0 1200 0 1 370
box -5 -3 28 105
use FILL  FILL_538
timestamp 1683038052
transform 1 0 1224 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1683038052
transform 1 0 1232 0 1 370
box -8 -3 104 105
use FILL  FILL_543
timestamp 1683038052
transform 1 0 1328 0 1 370
box -8 -3 16 105
use FILL  FILL_544
timestamp 1683038052
transform 1 0 1336 0 1 370
box -8 -3 16 105
use FILL  FILL_545
timestamp 1683038052
transform 1 0 1344 0 1 370
box -8 -3 16 105
use INVX2  INVX2_94
timestamp 1683038052
transform 1 0 1352 0 1 370
box -9 -3 26 105
use FILL  FILL_546
timestamp 1683038052
transform 1 0 1368 0 1 370
box -8 -3 16 105
use FILL  FILL_558
timestamp 1683038052
transform 1 0 1376 0 1 370
box -8 -3 16 105
use FILL  FILL_560
timestamp 1683038052
transform 1 0 1384 0 1 370
box -8 -3 16 105
use FILL  FILL_562
timestamp 1683038052
transform 1 0 1392 0 1 370
box -8 -3 16 105
use FILL  FILL_563
timestamp 1683038052
transform 1 0 1400 0 1 370
box -8 -3 16 105
use FILL  FILL_564
timestamp 1683038052
transform 1 0 1408 0 1 370
box -8 -3 16 105
use FILL  FILL_565
timestamp 1683038052
transform 1 0 1416 0 1 370
box -8 -3 16 105
use FILL  FILL_566
timestamp 1683038052
transform 1 0 1424 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_1014
timestamp 1683038052
transform 1 0 1444 0 1 375
box -3 -3 3 3
use INVX2  INVX2_96
timestamp 1683038052
transform 1 0 1432 0 1 370
box -9 -3 26 105
use FILL  FILL_567
timestamp 1683038052
transform 1 0 1448 0 1 370
box -8 -3 16 105
use FILL  FILL_568
timestamp 1683038052
transform 1 0 1456 0 1 370
box -8 -3 16 105
use FILL  FILL_569
timestamp 1683038052
transform 1 0 1464 0 1 370
box -8 -3 16 105
use FILL  FILL_570
timestamp 1683038052
transform 1 0 1472 0 1 370
box -8 -3 16 105
use FILL  FILL_571
timestamp 1683038052
transform 1 0 1480 0 1 370
box -8 -3 16 105
use FILL  FILL_572
timestamp 1683038052
transform 1 0 1488 0 1 370
box -8 -3 16 105
use FILL  FILL_573
timestamp 1683038052
transform 1 0 1496 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_1015
timestamp 1683038052
transform 1 0 1524 0 1 375
box -3 -3 3 3
use INVX2  INVX2_97
timestamp 1683038052
transform 1 0 1504 0 1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_51
timestamp 1683038052
transform 1 0 1520 0 1 370
box -8 -3 46 105
use FILL  FILL_574
timestamp 1683038052
transform 1 0 1560 0 1 370
box -8 -3 16 105
use FILL  FILL_575
timestamp 1683038052
transform 1 0 1568 0 1 370
box -8 -3 16 105
use INVX2  INVX2_98
timestamp 1683038052
transform 1 0 1576 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1683038052
transform 1 0 1592 0 1 370
box -8 -3 104 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_27
timestamp 1683038052
transform 1 0 1716 0 1 370
box -10 -3 10 3
use M2_M1  M2_M1_1201
timestamp 1683038052
transform 1 0 84 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1072
timestamp 1683038052
transform 1 0 84 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1683038052
transform 1 0 100 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1683038052
transform 1 0 116 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1683038052
transform 1 0 140 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1683038052
transform 1 0 132 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1683038052
transform 1 0 156 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1164
timestamp 1683038052
transform 1 0 100 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1683038052
transform 1 0 132 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1683038052
transform 1 0 140 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1683038052
transform 1 0 156 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1683038052
transform 1 0 172 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_1039
timestamp 1683038052
transform 1 0 180 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_1169
timestamp 1683038052
transform 1 0 196 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1170
timestamp 1683038052
transform 1 0 212 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1683038052
transform 1 0 228 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1683038052
transform 1 0 108 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1683038052
transform 1 0 124 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1683038052
transform 1 0 132 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1205
timestamp 1683038052
transform 1 0 148 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1048
timestamp 1683038052
transform 1 0 164 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_1206
timestamp 1683038052
transform 1 0 172 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1058
timestamp 1683038052
transform 1 0 132 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_1248
timestamp 1683038052
transform 1 0 172 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_1084
timestamp 1683038052
transform 1 0 108 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1073
timestamp 1683038052
transform 1 0 164 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1683038052
transform 1 0 252 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1683038052
transform 1 0 388 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_1156
timestamp 1683038052
transform 1 0 420 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1683038052
transform 1 0 316 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_1049
timestamp 1683038052
transform 1 0 212 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_1207
timestamp 1683038052
transform 1 0 252 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1050
timestamp 1683038052
transform 1 0 300 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1683038052
transform 1 0 420 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_1157
timestamp 1683038052
transform 1 0 444 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1683038052
transform 1 0 604 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1683038052
transform 1 0 428 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1683038052
transform 1 0 436 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1683038052
transform 1 0 548 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1208
timestamp 1683038052
transform 1 0 308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1209
timestamp 1683038052
transform 1 0 324 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1683038052
transform 1 0 332 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1042
timestamp 1683038052
transform 1 0 564 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1043
timestamp 1683038052
transform 1 0 580 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_1176
timestamp 1683038052
transform 1 0 604 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1683038052
transform 1 0 612 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1683038052
transform 1 0 532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1683038052
transform 1 0 540 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1051
timestamp 1683038052
transform 1 0 548 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_1213
timestamp 1683038052
transform 1 0 556 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1683038052
transform 1 0 564 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1215
timestamp 1683038052
transform 1 0 588 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1074
timestamp 1683038052
transform 1 0 196 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1683038052
transform 1 0 220 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1683038052
transform 1 0 308 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1683038052
transform 1 0 356 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1683038052
transform 1 0 412 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1683038052
transform 1 0 436 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1683038052
transform 1 0 508 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1683038052
transform 1 0 196 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1683038052
transform 1 0 292 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1683038052
transform 1 0 372 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1683038052
transform 1 0 404 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1683038052
transform 1 0 540 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1059
timestamp 1683038052
transform 1 0 604 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1683038052
transform 1 0 572 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1683038052
transform 1 0 612 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1683038052
transform 1 0 636 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1683038052
transform 1 0 708 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1683038052
transform 1 0 740 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_1178
timestamp 1683038052
transform 1 0 700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1683038052
transform 1 0 644 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1683038052
transform 1 0 652 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1218
timestamp 1683038052
transform 1 0 660 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1683038052
transform 1 0 684 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1029
timestamp 1683038052
transform 1 0 796 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1179
timestamp 1683038052
transform 1 0 756 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_1044
timestamp 1683038052
transform 1 0 764 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1683038052
transform 1 0 804 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_1220
timestamp 1683038052
transform 1 0 708 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1221
timestamp 1683038052
transform 1 0 716 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1222
timestamp 1683038052
transform 1 0 740 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1683038052
transform 1 0 756 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1683038052
transform 1 0 772 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1683038052
transform 1 0 796 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1683038052
transform 1 0 804 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1060
timestamp 1683038052
transform 1 0 660 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1683038052
transform 1 0 676 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1683038052
transform 1 0 700 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1063
timestamp 1683038052
transform 1 0 772 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_1180
timestamp 1683038052
transform 1 0 836 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1683038052
transform 1 0 852 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_1030
timestamp 1683038052
transform 1 0 860 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1181
timestamp 1683038052
transform 1 0 860 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_1046
timestamp 1683038052
transform 1 0 876 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1683038052
transform 1 0 908 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1683038052
transform 1 0 996 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1683038052
transform 1 0 900 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1032
timestamp 1683038052
transform 1 0 940 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1160
timestamp 1683038052
transform 1 0 1004 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1182
timestamp 1683038052
transform 1 0 884 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1683038052
transform 1 0 892 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1683038052
transform 1 0 900 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1683038052
transform 1 0 860 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1064
timestamp 1683038052
transform 1 0 860 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_1185
timestamp 1683038052
transform 1 0 1012 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1683038052
transform 1 0 1020 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1683038052
transform 1 0 892 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1683038052
transform 1 0 900 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1683038052
transform 1 0 916 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1065
timestamp 1683038052
transform 1 0 900 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1683038052
transform 1 0 1012 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1683038052
transform 1 0 1012 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1033
timestamp 1683038052
transform 1 0 1036 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1161
timestamp 1683038052
transform 1 0 1140 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1683038052
transform 1 0 1036 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1683038052
transform 1 0 1148 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1683038052
transform 1 0 1156 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1683038052
transform 1 0 1052 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1083
timestamp 1683038052
transform 1 0 1148 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1683038052
transform 1 0 1188 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1190
timestamp 1683038052
transform 1 0 1188 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1683038052
transform 1 0 1204 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1683038052
transform 1 0 1164 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1683038052
transform 1 0 1180 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1683038052
transform 1 0 1196 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1067
timestamp 1683038052
transform 1 0 1180 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1683038052
transform 1 0 1220 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_1235
timestamp 1683038052
transform 1 0 1228 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1683038052
transform 1 0 1244 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_1068
timestamp 1683038052
transform 1 0 1244 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1683038052
transform 1 0 1276 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_1236
timestamp 1683038052
transform 1 0 1268 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1683038052
transform 1 0 1276 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1683038052
transform 1 0 1292 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1035
timestamp 1683038052
transform 1 0 1348 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1194
timestamp 1683038052
transform 1 0 1332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1683038052
transform 1 0 1348 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_1053
timestamp 1683038052
transform 1 0 1332 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_1238
timestamp 1683038052
transform 1 0 1340 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1683038052
transform 1 0 1372 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_1054
timestamp 1683038052
transform 1 0 1372 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_1239
timestamp 1683038052
transform 1 0 1380 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1036
timestamp 1683038052
transform 1 0 1420 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1197
timestamp 1683038052
transform 1 0 1404 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1683038052
transform 1 0 1420 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_1026
timestamp 1683038052
transform 1 0 1548 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_1162
timestamp 1683038052
transform 1 0 1444 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_1037
timestamp 1683038052
transform 1 0 1548 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1683038052
transform 1 0 1540 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_1199
timestamp 1683038052
transform 1 0 1548 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1683038052
transform 1 0 1396 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1241
timestamp 1683038052
transform 1 0 1412 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1683038052
transform 1 0 1428 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1055
timestamp 1683038052
transform 1 0 1508 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_1243
timestamp 1683038052
transform 1 0 1532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1244
timestamp 1683038052
transform 1 0 1540 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1056
timestamp 1683038052
transform 1 0 1548 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1069
timestamp 1683038052
transform 1 0 1540 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_1163
timestamp 1683038052
transform 1 0 1580 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_1038
timestamp 1683038052
transform 1 0 1692 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1200
timestamp 1683038052
transform 1 0 1692 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1683038052
transform 1 0 1564 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1057
timestamp 1683038052
transform 1 0 1572 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_1246
timestamp 1683038052
transform 1 0 1668 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1683038052
transform 1 0 1676 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1070
timestamp 1683038052
transform 1 0 1564 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1071
timestamp 1683038052
transform 1 0 1676 0 1 315
box -3 -3 3 3
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_28
timestamp 1683038052
transform 1 0 24 0 1 270
box -10 -3 10 3
use M3_M2  M3_M2_1091
timestamp 1683038052
transform 1 0 68 0 1 275
box -3 -3 3 3
use FILL  FILL_508
timestamp 1683038052
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_509
timestamp 1683038052
transform 1 0 80 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_46
timestamp 1683038052
transform 1 0 88 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_47
timestamp 1683038052
transform 1 0 128 0 -1 370
box -8 -3 46 105
use M3_M2  M3_M2_1092
timestamp 1683038052
transform 1 0 180 0 1 275
box -3 -3 3 3
use OAI21X1  OAI21X1_36
timestamp 1683038052
transform -1 0 200 0 -1 370
box -8 -3 34 105
use INVX2  INVX2_88
timestamp 1683038052
transform -1 0 216 0 -1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1683038052
transform 1 0 216 0 -1 370
box -8 -3 104 105
use FAX1  FAX1_21
timestamp 1683038052
transform 1 0 312 0 -1 370
box -5 -3 126 105
use FAX1  FAX1_22
timestamp 1683038052
transform -1 0 552 0 -1 370
box -5 -3 126 105
use MUX2X1  MUX2X1_18
timestamp 1683038052
transform 1 0 552 0 -1 370
box -5 -3 53 105
use NOR2X1  NOR2X1_17
timestamp 1683038052
transform 1 0 600 0 -1 370
box -8 -3 32 105
use FILL  FILL_517
timestamp 1683038052
transform 1 0 624 0 -1 370
box -8 -3 16 105
use FILL  FILL_518
timestamp 1683038052
transform 1 0 632 0 -1 370
box -8 -3 16 105
use FILL  FILL_519
timestamp 1683038052
transform 1 0 640 0 -1 370
box -8 -3 16 105
use MUX2X1  MUX2X1_21
timestamp 1683038052
transform 1 0 648 0 -1 370
box -5 -3 53 105
use FILL  FILL_520
timestamp 1683038052
transform 1 0 696 0 -1 370
box -8 -3 16 105
use MUX2X1  MUX2X1_22
timestamp 1683038052
transform 1 0 704 0 -1 370
box -5 -3 53 105
use FILL  FILL_521
timestamp 1683038052
transform 1 0 752 0 -1 370
box -8 -3 16 105
use MUX2X1  MUX2X1_23
timestamp 1683038052
transform 1 0 760 0 -1 370
box -5 -3 53 105
use FILL  FILL_522
timestamp 1683038052
transform 1 0 808 0 -1 370
box -8 -3 16 105
use FILL  FILL_523
timestamp 1683038052
transform 1 0 816 0 -1 370
box -8 -3 16 105
use FILL  FILL_539
timestamp 1683038052
transform 1 0 824 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_18
timestamp 1683038052
transform -1 0 856 0 -1 370
box -8 -3 32 105
use INVX2  INVX2_91
timestamp 1683038052
transform 1 0 856 0 -1 370
box -9 -3 26 105
use NOR2X1  NOR2X1_19
timestamp 1683038052
transform 1 0 872 0 -1 370
box -8 -3 32 105
use FAX1  FAX1_23
timestamp 1683038052
transform 1 0 896 0 -1 370
box -5 -3 126 105
use INVX2  INVX2_92
timestamp 1683038052
transform 1 0 1016 0 -1 370
box -9 -3 26 105
use M3_M2  M3_M2_1093
timestamp 1683038052
transform 1 0 1148 0 1 275
box -3 -3 3 3
use FAX1  FAX1_24
timestamp 1683038052
transform 1 0 1032 0 -1 370
box -5 -3 126 105
use FILL  FILL_540
timestamp 1683038052
transform 1 0 1152 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_1094
timestamp 1683038052
transform 1 0 1204 0 1 275
box -3 -3 3 3
use AOI22X1  AOI22X1_49
timestamp 1683038052
transform 1 0 1160 0 -1 370
box -8 -3 46 105
use INVX2  INVX2_93
timestamp 1683038052
transform 1 0 1200 0 -1 370
box -9 -3 26 105
use FILL  FILL_541
timestamp 1683038052
transform 1 0 1216 0 -1 370
box -8 -3 16 105
use FILL  FILL_542
timestamp 1683038052
transform 1 0 1224 0 -1 370
box -8 -3 16 105
use FILL  FILL_547
timestamp 1683038052
transform 1 0 1232 0 -1 370
box -8 -3 16 105
use FILL  FILL_548
timestamp 1683038052
transform 1 0 1240 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_95
timestamp 1683038052
transform 1 0 1248 0 -1 370
box -9 -3 26 105
use FILL  FILL_549
timestamp 1683038052
transform 1 0 1264 0 -1 370
box -8 -3 16 105
use FILL  FILL_550
timestamp 1683038052
transform 1 0 1272 0 -1 370
box -8 -3 16 105
use FILL  FILL_551
timestamp 1683038052
transform 1 0 1280 0 -1 370
box -8 -3 16 105
use FILL  FILL_552
timestamp 1683038052
transform 1 0 1288 0 -1 370
box -8 -3 16 105
use FILL  FILL_553
timestamp 1683038052
transform 1 0 1296 0 -1 370
box -8 -3 16 105
use FILL  FILL_554
timestamp 1683038052
transform 1 0 1304 0 -1 370
box -8 -3 16 105
use FILL  FILL_555
timestamp 1683038052
transform 1 0 1312 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_50
timestamp 1683038052
transform 1 0 1320 0 -1 370
box -8 -3 46 105
use FILL  FILL_556
timestamp 1683038052
transform 1 0 1360 0 -1 370
box -8 -3 16 105
use FILL  FILL_557
timestamp 1683038052
transform 1 0 1368 0 -1 370
box -8 -3 16 105
use FILL  FILL_559
timestamp 1683038052
transform 1 0 1376 0 -1 370
box -8 -3 16 105
use FILL  FILL_561
timestamp 1683038052
transform 1 0 1384 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_52
timestamp 1683038052
transform 1 0 1392 0 -1 370
box -8 -3 46 105
use FAX1  FAX1_25
timestamp 1683038052
transform -1 0 1552 0 -1 370
box -5 -3 126 105
use INVX2  INVX2_99
timestamp 1683038052
transform 1 0 1552 0 -1 370
box -9 -3 26 105
use FAX1  FAX1_26
timestamp 1683038052
transform -1 0 1688 0 -1 370
box -5 -3 126 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_29
timestamp 1683038052
transform 1 0 1740 0 1 270
box -10 -3 10 3
use M3_M2  M3_M2_1114
timestamp 1683038052
transform 1 0 84 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1115
timestamp 1683038052
transform 1 0 124 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1116
timestamp 1683038052
transform 1 0 140 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1117
timestamp 1683038052
transform 1 0 180 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1250
timestamp 1683038052
transform 1 0 68 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1683038052
transform 1 0 140 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1683038052
transform 1 0 180 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1683038052
transform 1 0 164 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1683038052
transform 1 0 196 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1683038052
transform 1 0 188 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1683038052
transform 1 0 196 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1161
timestamp 1683038052
transform 1 0 188 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_1297
timestamp 1683038052
transform 1 0 220 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1095
timestamp 1683038052
transform 1 0 244 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1096
timestamp 1683038052
transform 1 0 332 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_1253
timestamp 1683038052
transform 1 0 340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1683038052
transform 1 0 236 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1299
timestamp 1683038052
transform 1 0 244 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1149
timestamp 1683038052
transform 1 0 252 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_1300
timestamp 1683038052
transform 1 0 356 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1683038052
transform 1 0 252 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1683038052
transform 1 0 380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1683038052
transform 1 0 396 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1132
timestamp 1683038052
transform 1 0 404 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1256
timestamp 1683038052
transform 1 0 412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1257
timestamp 1683038052
transform 1 0 420 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1683038052
transform 1 0 436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1683038052
transform 1 0 372 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1150
timestamp 1683038052
transform 1 0 380 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1683038052
transform 1 0 444 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1302
timestamp 1683038052
transform 1 0 388 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1683038052
transform 1 0 404 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1683038052
transform 1 0 412 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1683038052
transform 1 0 428 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1683038052
transform 1 0 444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1683038052
transform 1 0 452 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1169
timestamp 1683038052
transform 1 0 236 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1170
timestamp 1683038052
transform 1 0 284 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1683038052
transform 1 0 364 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1683038052
transform 1 0 396 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1172
timestamp 1683038052
transform 1 0 452 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1683038052
transform 1 0 556 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1683038052
transform 1 0 588 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1118
timestamp 1683038052
transform 1 0 564 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1683038052
transform 1 0 636 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1683038052
transform 1 0 700 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1259
timestamp 1683038052
transform 1 0 524 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1683038052
transform 1 0 540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1683038052
transform 1 0 548 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1683038052
transform 1 0 556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1683038052
transform 1 0 588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1264
timestamp 1683038052
transform 1 0 596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1683038052
transform 1 0 604 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1683038052
transform 1 0 636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1683038052
transform 1 0 644 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1683038052
transform 1 0 652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1683038052
transform 1 0 676 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1683038052
transform 1 0 508 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1151
timestamp 1683038052
transform 1 0 548 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1152
timestamp 1683038052
transform 1 0 572 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_1309
timestamp 1683038052
transform 1 0 588 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1153
timestamp 1683038052
transform 1 0 596 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1154
timestamp 1683038052
transform 1 0 620 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_1310
timestamp 1683038052
transform 1 0 636 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1173
timestamp 1683038052
transform 1 0 524 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1683038052
transform 1 0 596 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1683038052
transform 1 0 692 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1270
timestamp 1683038052
transform 1 0 700 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1683038052
transform 1 0 708 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1135
timestamp 1683038052
transform 1 0 716 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1272
timestamp 1683038052
transform 1 0 732 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1136
timestamp 1683038052
transform 1 0 740 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1311
timestamp 1683038052
transform 1 0 692 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1155
timestamp 1683038052
transform 1 0 740 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1121
timestamp 1683038052
transform 1 0 756 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1683038052
transform 1 0 796 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1273
timestamp 1683038052
transform 1 0 756 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1683038052
transform 1 0 764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1683038052
transform 1 0 788 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1683038052
transform 1 0 748 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1175
timestamp 1683038052
transform 1 0 708 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1683038052
transform 1 0 804 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1313
timestamp 1683038052
transform 1 0 796 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1683038052
transform 1 0 804 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1683038052
transform 1 0 844 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1683038052
transform 1 0 852 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1156
timestamp 1683038052
transform 1 0 844 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1683038052
transform 1 0 868 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1315
timestamp 1683038052
transform 1 0 860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1683038052
transform 1 0 868 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1157
timestamp 1683038052
transform 1 0 876 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1163
timestamp 1683038052
transform 1 0 860 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_1337
timestamp 1683038052
transform 1 0 876 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_1123
timestamp 1683038052
transform 1 0 900 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1278
timestamp 1683038052
transform 1 0 892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1683038052
transform 1 0 900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1683038052
transform 1 0 900 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1139
timestamp 1683038052
transform 1 0 916 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1338
timestamp 1683038052
transform 1 0 916 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_1176
timestamp 1683038052
transform 1 0 908 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1683038052
transform 1 0 940 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1683038052
transform 1 0 956 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_1318
timestamp 1683038052
transform 1 0 948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1683038052
transform 1 0 972 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1178
timestamp 1683038052
transform 1 0 972 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1107
timestamp 1683038052
transform 1 0 1028 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1108
timestamp 1683038052
transform 1 0 1044 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_1280
timestamp 1683038052
transform 1 0 1012 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1140
timestamp 1683038052
transform 1 0 1044 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1141
timestamp 1683038052
transform 1 0 1108 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1158
timestamp 1683038052
transform 1 0 1100 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_1320
timestamp 1683038052
transform 1 0 1108 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1683038052
transform 1 0 1116 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1097
timestamp 1683038052
transform 1 0 1156 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1683038052
transform 1 0 1188 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1099
timestamp 1683038052
transform 1 0 1196 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1683038052
transform 1 0 1164 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1124
timestamp 1683038052
transform 1 0 1124 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1683038052
transform 1 0 1348 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1111
timestamp 1683038052
transform 1 0 1364 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1112
timestamp 1683038052
transform 1 0 1380 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1100
timestamp 1683038052
transform 1 0 1420 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1683038052
transform 1 0 1428 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1683038052
transform 1 0 1556 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1125
timestamp 1683038052
transform 1 0 1172 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1683038052
transform 1 0 1284 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1127
timestamp 1683038052
transform 1 0 1308 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1683038052
transform 1 0 1404 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1683038052
transform 1 0 1428 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1130
timestamp 1683038052
transform 1 0 1524 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1281
timestamp 1683038052
transform 1 0 1124 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1683038052
transform 1 0 1132 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1683038052
transform 1 0 1148 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1683038052
transform 1 0 1164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1285
timestamp 1683038052
transform 1 0 1172 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1164
timestamp 1683038052
transform 1 0 1076 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_1339
timestamp 1683038052
transform 1 0 1100 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_1165
timestamp 1683038052
transform 1 0 1116 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1683038052
transform 1 0 1044 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1683038052
transform 1 0 1180 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1286
timestamp 1683038052
transform 1 0 1188 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1143
timestamp 1683038052
transform 1 0 1276 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1144
timestamp 1683038052
transform 1 0 1292 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1287
timestamp 1683038052
transform 1 0 1300 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1288
timestamp 1683038052
transform 1 0 1308 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1145
timestamp 1683038052
transform 1 0 1396 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1146
timestamp 1683038052
transform 1 0 1412 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1289
timestamp 1683038052
transform 1 0 1420 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1683038052
transform 1 0 1428 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1147
timestamp 1683038052
transform 1 0 1444 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1683038052
transform 1 0 1532 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1291
timestamp 1683038052
transform 1 0 1548 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1683038052
transform 1 0 1140 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1683038052
transform 1 0 1156 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1159
timestamp 1683038052
transform 1 0 1164 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_1324
timestamp 1683038052
transform 1 0 1172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1683038052
transform 1 0 1284 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1683038052
transform 1 0 1292 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1180
timestamp 1683038052
transform 1 0 1132 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1160
timestamp 1683038052
transform 1 0 1308 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_1327
timestamp 1683038052
transform 1 0 1404 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1683038052
transform 1 0 1412 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1166
timestamp 1683038052
transform 1 0 1172 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_1340
timestamp 1683038052
transform 1 0 1276 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_1167
timestamp 1683038052
transform 1 0 1292 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_1341
timestamp 1683038052
transform 1 0 1396 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_1102
timestamp 1683038052
transform 1 0 1580 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1683038052
transform 1 0 1684 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1683038052
transform 1 0 1588 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1292
timestamp 1683038052
transform 1 0 1580 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1683038052
transform 1 0 1588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1683038052
transform 1 0 1524 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1683038052
transform 1 0 1532 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1683038052
transform 1 0 1540 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1683038052
transform 1 0 1556 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1333
timestamp 1683038052
transform 1 0 1564 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1683038052
transform 1 0 1572 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1683038052
transform 1 0 1692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1683038052
transform 1 0 1516 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_1181
timestamp 1683038052
transform 1 0 1516 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1683038052
transform 1 0 1572 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_1343
timestamp 1683038052
transform 1 0 1676 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_1182
timestamp 1683038052
transform 1 0 1564 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1183
timestamp 1683038052
transform 1 0 1676 0 1 185
box -3 -3 3 3
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_30
timestamp 1683038052
transform 1 0 48 0 1 170
box -10 -3 10 3
use FILL  FILL_576
timestamp 1683038052
transform 1 0 72 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1683038052
transform -1 0 176 0 1 170
box -8 -3 104 105
use INVX2  INVX2_100
timestamp 1683038052
transform -1 0 192 0 1 170
box -9 -3 26 105
use OAI21X1  OAI21X1_37
timestamp 1683038052
transform -1 0 224 0 1 170
box -8 -3 34 105
use INVX2  INVX2_101
timestamp 1683038052
transform -1 0 240 0 1 170
box -9 -3 26 105
use FAX1  FAX1_27
timestamp 1683038052
transform -1 0 360 0 1 170
box -5 -3 126 105
use INVX2  INVX2_102
timestamp 1683038052
transform -1 0 376 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_53
timestamp 1683038052
transform 1 0 376 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_54
timestamp 1683038052
transform 1 0 416 0 1 170
box -8 -3 46 105
use XOR2X1  XOR2X1_5
timestamp 1683038052
transform -1 0 512 0 1 170
box -8 -3 64 105
use AND2X2  AND2X2_6
timestamp 1683038052
transform 1 0 512 0 1 170
box -8 -3 40 105
use MUX2X1  MUX2X1_25
timestamp 1683038052
transform 1 0 544 0 1 170
box -5 -3 53 105
use MUX2X1  MUX2X1_26
timestamp 1683038052
transform 1 0 592 0 1 170
box -5 -3 53 105
use MUX2X1  MUX2X1_27
timestamp 1683038052
transform 1 0 640 0 1 170
box -5 -3 53 105
use FILL  FILL_578
timestamp 1683038052
transform 1 0 688 0 1 170
box -8 -3 16 105
use MUX2X1  MUX2X1_28
timestamp 1683038052
transform 1 0 696 0 1 170
box -5 -3 53 105
use FILL  FILL_579
timestamp 1683038052
transform 1 0 744 0 1 170
box -8 -3 16 105
use MUX2X1  MUX2X1_29
timestamp 1683038052
transform 1 0 752 0 1 170
box -5 -3 53 105
use INVX2  INVX2_103
timestamp 1683038052
transform 1 0 800 0 1 170
box -9 -3 26 105
use FILL  FILL_604
timestamp 1683038052
transform 1 0 816 0 1 170
box -8 -3 16 105
use FILL  FILL_605
timestamp 1683038052
transform 1 0 824 0 1 170
box -8 -3 16 105
use FILL  FILL_606
timestamp 1683038052
transform 1 0 832 0 1 170
box -8 -3 16 105
use FILL  FILL_608
timestamp 1683038052
transform 1 0 840 0 1 170
box -8 -3 16 105
use NOR2X1  NOR2X1_21
timestamp 1683038052
transform -1 0 872 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_22
timestamp 1683038052
transform 1 0 872 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_23
timestamp 1683038052
transform -1 0 920 0 1 170
box -8 -3 32 105
use FILL  FILL_609
timestamp 1683038052
transform 1 0 920 0 1 170
box -8 -3 16 105
use FILL  FILL_615
timestamp 1683038052
transform 1 0 928 0 1 170
box -8 -3 16 105
use FILL  FILL_617
timestamp 1683038052
transform 1 0 936 0 1 170
box -8 -3 16 105
use FILL  FILL_618
timestamp 1683038052
transform 1 0 944 0 1 170
box -8 -3 16 105
use INVX2  INVX2_108
timestamp 1683038052
transform 1 0 952 0 1 170
box -9 -3 26 105
use FILL  FILL_619
timestamp 1683038052
transform 1 0 968 0 1 170
box -8 -3 16 105
use FILL  FILL_620
timestamp 1683038052
transform 1 0 976 0 1 170
box -8 -3 16 105
use FILL  FILL_621
timestamp 1683038052
transform 1 0 984 0 1 170
box -8 -3 16 105
use FAX1  FAX1_28
timestamp 1683038052
transform 1 0 992 0 1 170
box -5 -3 126 105
use INVX2  INVX2_109
timestamp 1683038052
transform 1 0 1112 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_55
timestamp 1683038052
transform 1 0 1128 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_1184
timestamp 1683038052
transform 1 0 1196 0 1 175
box -3 -3 3 3
use FAX1  FAX1_29
timestamp 1683038052
transform 1 0 1168 0 1 170
box -5 -3 126 105
use M3_M2  M3_M2_1185
timestamp 1683038052
transform 1 0 1300 0 1 175
box -3 -3 3 3
use FAX1  FAX1_30
timestamp 1683038052
transform 1 0 1288 0 1 170
box -5 -3 126 105
use FAX1  FAX1_31
timestamp 1683038052
transform 1 0 1408 0 1 170
box -5 -3 126 105
use AOI22X1  AOI22X1_56
timestamp 1683038052
transform 1 0 1528 0 1 170
box -8 -3 46 105
use FAX1  FAX1_32
timestamp 1683038052
transform 1 0 1568 0 1 170
box -5 -3 126 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_31
timestamp 1683038052
transform 1 0 1716 0 1 170
box -10 -3 10 3
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_32
timestamp 1683038052
transform 1 0 24 0 1 70
box -10 -3 10 3
use M2_M1  M2_M1_1353
timestamp 1683038052
transform 1 0 164 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1683038052
transform 1 0 84 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1683038052
transform 1 0 140 0 1 125
box -2 -2 2 2
use FILL  FILL_577
timestamp 1683038052
transform 1 0 72 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1226
timestamp 1683038052
transform 1 0 140 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_64
timestamp 1683038052
transform -1 0 176 0 -1 170
box -8 -3 104 105
use FILL  FILL_580
timestamp 1683038052
transform 1 0 176 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1186
timestamp 1683038052
transform 1 0 204 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1683038052
transform 1 0 228 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1683038052
transform 1 0 196 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1683038052
transform 1 0 228 0 1 155
box -3 -3 3 3
use FILL  FILL_581
timestamp 1683038052
transform 1 0 184 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1354
timestamp 1683038052
transform 1 0 204 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1683038052
transform 1 0 228 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1683038052
transform 1 0 284 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1683038052
transform 1 0 292 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1227
timestamp 1683038052
transform 1 0 292 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_65
timestamp 1683038052
transform 1 0 192 0 -1 170
box -8 -3 104 105
use FILL  FILL_582
timestamp 1683038052
transform 1 0 288 0 -1 170
box -8 -3 16 105
use FILL  FILL_583
timestamp 1683038052
transform 1 0 296 0 -1 170
box -8 -3 16 105
use INVX2  INVX2_104
timestamp 1683038052
transform -1 0 320 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_1188
timestamp 1683038052
transform 1 0 332 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_1355
timestamp 1683038052
transform 1 0 332 0 1 135
box -2 -2 2 2
use FILL  FILL_584
timestamp 1683038052
transform 1 0 320 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1384
timestamp 1683038052
transform 1 0 340 0 1 125
box -2 -2 2 2
use FILL  FILL_585
timestamp 1683038052
transform 1 0 328 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1344
timestamp 1683038052
transform 1 0 364 0 1 145
box -2 -2 2 2
use OR2X1  OR2X1_4
timestamp 1683038052
transform -1 0 368 0 -1 170
box -8 -3 40 105
use FILL  FILL_586
timestamp 1683038052
transform 1 0 368 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1195
timestamp 1683038052
transform 1 0 396 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1683038052
transform 1 0 388 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1356
timestamp 1683038052
transform 1 0 388 0 1 135
box -2 -2 2 2
use FILL  FILL_587
timestamp 1683038052
transform 1 0 376 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1385
timestamp 1683038052
transform 1 0 396 0 1 125
box -2 -2 2 2
use FILL  FILL_588
timestamp 1683038052
transform 1 0 384 0 -1 170
box -8 -3 16 105
use FILL  FILL_589
timestamp 1683038052
transform 1 0 392 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1189
timestamp 1683038052
transform 1 0 436 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1683038052
transform 1 0 420 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1209
timestamp 1683038052
transform 1 0 452 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1357
timestamp 1683038052
transform 1 0 452 0 1 135
box -2 -2 2 2
use XNOR2X1  XNOR2X1_4
timestamp 1683038052
transform -1 0 456 0 -1 170
box -8 -3 64 105
use FILL  FILL_590
timestamp 1683038052
transform 1 0 456 0 -1 170
box -8 -3 16 105
use FILL  FILL_591
timestamp 1683038052
transform 1 0 464 0 -1 170
box -8 -3 16 105
use FILL  FILL_592
timestamp 1683038052
transform 1 0 472 0 -1 170
box -8 -3 16 105
use FILL  FILL_593
timestamp 1683038052
transform 1 0 480 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1358
timestamp 1683038052
transform 1 0 508 0 1 135
box -2 -2 2 2
use INVX2  INVX2_105
timestamp 1683038052
transform -1 0 504 0 -1 170
box -9 -3 26 105
use FILL  FILL_594
timestamp 1683038052
transform 1 0 504 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1386
timestamp 1683038052
transform 1 0 524 0 1 125
box -2 -2 2 2
use FILL  FILL_595
timestamp 1683038052
transform 1 0 512 0 -1 170
box -8 -3 16 105
use FILL  FILL_596
timestamp 1683038052
transform 1 0 520 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1359
timestamp 1683038052
transform 1 0 540 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_1219
timestamp 1683038052
transform 1 0 548 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_1387
timestamp 1683038052
transform 1 0 564 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1683038052
transform 1 0 572 0 1 125
box -2 -2 2 2
use MUX2X1  MUX2X1_30
timestamp 1683038052
transform -1 0 576 0 -1 170
box -5 -3 53 105
use M2_M1  M2_M1_1360
timestamp 1683038052
transform 1 0 596 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_1220
timestamp 1683038052
transform 1 0 620 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1683038052
transform 1 0 684 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1210
timestamp 1683038052
transform 1 0 724 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1345
timestamp 1683038052
transform 1 0 740 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1683038052
transform 1 0 684 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1683038052
transform 1 0 724 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1683038052
transform 1 0 588 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1683038052
transform 1 0 620 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1683038052
transform 1 0 636 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1683038052
transform 1 0 644 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1683038052
transform 1 0 668 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1683038052
transform 1 0 676 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1228
timestamp 1683038052
transform 1 0 588 0 1 115
box -3 -3 3 3
use FILL  FILL_597
timestamp 1683038052
transform 1 0 576 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1229
timestamp 1683038052
transform 1 0 644 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1683038052
transform 1 0 668 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1240
timestamp 1683038052
transform 1 0 636 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1241
timestamp 1683038052
transform 1 0 660 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1683038052
transform 1 0 676 0 1 105
box -3 -3 3 3
use MUX2X1  MUX2X1_31
timestamp 1683038052
transform -1 0 632 0 -1 170
box -5 -3 53 105
use MUX2X1  MUX2X1_32
timestamp 1683038052
transform 1 0 632 0 -1 170
box -5 -3 53 105
use FILL  FILL_598
timestamp 1683038052
transform 1 0 680 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1198
timestamp 1683038052
transform 1 0 764 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1395
timestamp 1683038052
transform 1 0 700 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1683038052
transform 1 0 740 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1683038052
transform 1 0 756 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1231
timestamp 1683038052
transform 1 0 700 0 1 115
box -3 -3 3 3
use MUX2X1  MUX2X1_33
timestamp 1683038052
transform 1 0 688 0 -1 170
box -5 -3 53 105
use M3_M2  M3_M2_1243
timestamp 1683038052
transform 1 0 756 0 1 105
box -3 -3 3 3
use NOR2X1  NOR2X1_20
timestamp 1683038052
transform 1 0 736 0 -1 170
box -8 -3 32 105
use FILL  FILL_599
timestamp 1683038052
transform 1 0 760 0 -1 170
box -8 -3 16 105
use FILL  FILL_600
timestamp 1683038052
transform 1 0 768 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1346
timestamp 1683038052
transform 1 0 788 0 1 145
box -2 -2 2 2
use FILL  FILL_601
timestamp 1683038052
transform 1 0 776 0 -1 170
box -8 -3 16 105
use FILL  FILL_602
timestamp 1683038052
transform 1 0 784 0 -1 170
box -8 -3 16 105
use FILL  FILL_603
timestamp 1683038052
transform 1 0 792 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1211
timestamp 1683038052
transform 1 0 820 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1683038052
transform 1 0 812 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_1363
timestamp 1683038052
transform 1 0 820 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1683038052
transform 1 0 812 0 1 125
box -2 -2 2 2
use INVX2  INVX2_106
timestamp 1683038052
transform 1 0 800 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_107
timestamp 1683038052
transform 1 0 816 0 -1 170
box -9 -3 26 105
use FILL  FILL_607
timestamp 1683038052
transform 1 0 832 0 -1 170
box -8 -3 16 105
use FILL  FILL_610
timestamp 1683038052
transform 1 0 840 0 -1 170
box -8 -3 16 105
use FILL  FILL_611
timestamp 1683038052
transform 1 0 848 0 -1 170
box -8 -3 16 105
use FILL  FILL_612
timestamp 1683038052
transform 1 0 856 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1190
timestamp 1683038052
transform 1 0 900 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1212
timestamp 1683038052
transform 1 0 892 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1364
timestamp 1683038052
transform 1 0 892 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1683038052
transform 1 0 884 0 1 125
box -2 -2 2 2
use NOR2X1  NOR2X1_24
timestamp 1683038052
transform 1 0 864 0 -1 170
box -8 -3 32 105
use M2_M1  M2_M1_1347
timestamp 1683038052
transform 1 0 908 0 1 145
box -2 -2 2 2
use M3_M2  M3_M2_1222
timestamp 1683038052
transform 1 0 908 0 1 135
box -3 -3 3 3
use NOR2X1  NOR2X1_25
timestamp 1683038052
transform -1 0 912 0 -1 170
box -8 -3 32 105
use FILL  FILL_613
timestamp 1683038052
transform 1 0 912 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1199
timestamp 1683038052
transform 1 0 1052 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1348
timestamp 1683038052
transform 1 0 1044 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1365
timestamp 1683038052
transform 1 0 932 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1366
timestamp 1683038052
transform 1 0 940 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_1223
timestamp 1683038052
transform 1 0 932 0 1 125
box -3 -3 3 3
use FILL  FILL_614
timestamp 1683038052
transform 1 0 920 0 -1 170
box -8 -3 16 105
use FILL  FILL_616
timestamp 1683038052
transform 1 0 928 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1200
timestamp 1683038052
transform 1 0 1068 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1683038052
transform 1 0 1180 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1191
timestamp 1683038052
transform 1 0 1324 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1683038052
transform 1 0 1348 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1683038052
transform 1 0 1204 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1203
timestamp 1683038052
transform 1 0 1292 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1349
timestamp 1683038052
transform 1 0 1172 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1683038052
transform 1 0 1060 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1683038052
transform 1 0 1068 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1400
timestamp 1683038052
transform 1 0 948 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1401
timestamp 1683038052
transform 1 0 956 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1213
timestamp 1683038052
transform 1 0 1188 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1683038052
transform 1 0 1212 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1350
timestamp 1683038052
transform 1 0 1308 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1683038052
transform 1 0 1180 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1370
timestamp 1683038052
transform 1 0 1188 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1683038052
transform 1 0 1076 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1683038052
transform 1 0 1084 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1683038052
transform 1 0 1204 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_1204
timestamp 1683038052
transform 1 0 1340 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1683038052
transform 1 0 1412 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1683038052
transform 1 0 1532 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1683038052
transform 1 0 1564 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1683038052
transform 1 0 1332 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1683038052
transform 1 0 1420 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1351
timestamp 1683038052
transform 1 0 1444 0 1 145
box -2 -2 2 2
use M3_M2  M3_M2_1217
timestamp 1683038052
transform 1 0 1460 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1352
timestamp 1683038052
transform 1 0 1564 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1683038052
transform 1 0 1316 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1683038052
transform 1 0 1324 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1683038052
transform 1 0 1196 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1683038052
transform 1 0 1212 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1683038052
transform 1 0 1220 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1232
timestamp 1683038052
transform 1 0 1060 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1683038052
transform 1 0 1084 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1683038052
transform 1 0 1180 0 1 115
box -3 -3 3 3
use FAX1  FAX1_33
timestamp 1683038052
transform 1 0 936 0 -1 170
box -5 -3 126 105
use FILL  FILL_622
timestamp 1683038052
transform 1 0 1056 0 -1 170
box -8 -3 16 105
use FAX1  FAX1_34
timestamp 1683038052
transform 1 0 1064 0 -1 170
box -5 -3 126 105
use INVX2  INVX2_110
timestamp 1683038052
transform 1 0 1184 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_1374
timestamp 1683038052
transform 1 0 1340 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1683038052
transform 1 0 1452 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1376
timestamp 1683038052
transform 1 0 1460 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_1218
timestamp 1683038052
transform 1 0 1580 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1377
timestamp 1683038052
transform 1 0 1572 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1683038052
transform 1 0 1332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1683038052
transform 1 0 1348 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1683038052
transform 1 0 1356 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1235
timestamp 1683038052
transform 1 0 1220 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1683038052
transform 1 0 1316 0 1 115
box -3 -3 3 3
use FAX1  FAX1_35
timestamp 1683038052
transform 1 0 1200 0 -1 170
box -5 -3 126 105
use INVX2  INVX2_111
timestamp 1683038052
transform 1 0 1320 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_1224
timestamp 1683038052
transform 1 0 1452 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_1410
timestamp 1683038052
transform 1 0 1460 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1225
timestamp 1683038052
transform 1 0 1468 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_1411
timestamp 1683038052
transform 1 0 1476 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1237
timestamp 1683038052
transform 1 0 1356 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1683038052
transform 1 0 1460 0 1 115
box -3 -3 3 3
use FAX1  FAX1_36
timestamp 1683038052
transform 1 0 1336 0 -1 170
box -5 -3 126 105
use FAX1  FAX1_37
timestamp 1683038052
transform 1 0 1456 0 -1 170
box -5 -3 126 105
use M2_M1  M2_M1_1378
timestamp 1683038052
transform 1 0 1588 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_1239
timestamp 1683038052
transform 1 0 1588 0 1 115
box -3 -3 3 3
use FILL  FILL_623
timestamp 1683038052
transform 1 0 1576 0 -1 170
box -8 -3 16 105
use FILL  FILL_624
timestamp 1683038052
transform 1 0 1584 0 -1 170
box -8 -3 16 105
use INVX2  INVX2_112
timestamp 1683038052
transform 1 0 1592 0 -1 170
box -9 -3 26 105
use FILL  FILL_625
timestamp 1683038052
transform 1 0 1608 0 -1 170
box -8 -3 16 105
use FILL  FILL_626
timestamp 1683038052
transform 1 0 1616 0 -1 170
box -8 -3 16 105
use FILL  FILL_627
timestamp 1683038052
transform 1 0 1624 0 -1 170
box -8 -3 16 105
use FILL  FILL_628
timestamp 1683038052
transform 1 0 1632 0 -1 170
box -8 -3 16 105
use FILL  FILL_629
timestamp 1683038052
transform 1 0 1640 0 -1 170
box -8 -3 16 105
use FILL  FILL_630
timestamp 1683038052
transform 1 0 1648 0 -1 170
box -8 -3 16 105
use FILL  FILL_631
timestamp 1683038052
transform 1 0 1656 0 -1 170
box -8 -3 16 105
use FILL  FILL_632
timestamp 1683038052
transform 1 0 1664 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1412
timestamp 1683038052
transform 1 0 1684 0 1 125
box -2 -2 2 2
use FILL  FILL_633
timestamp 1683038052
transform 1 0 1672 0 -1 170
box -8 -3 16 105
use FILL  FILL_634
timestamp 1683038052
transform 1 0 1680 0 -1 170
box -8 -3 16 105
use CORDIC_TOP_VIA0  CORDIC_TOP_VIA0_33
timestamp 1683038052
transform 1 0 1740 0 1 70
box -10 -3 10 3
use CORDIC_TOP_VIA1  CORDIC_TOP_VIA1_4
timestamp 1683038052
transform 1 0 48 0 1 47
box -10 -10 10 10
use CORDIC_TOP_VIA1  CORDIC_TOP_VIA1_5
timestamp 1683038052
transform 1 0 1716 0 1 47
box -10 -10 10 10
use CORDIC_TOP_VIA1  CORDIC_TOP_VIA1_6
timestamp 1683038052
transform 1 0 24 0 1 23
box -10 -10 10 10
use CORDIC_TOP_VIA1  CORDIC_TOP_VIA1_7
timestamp 1683038052
transform 1 0 1740 0 1 23
box -10 -10 10 10
<< labels >>
rlabel metal2 860 1738 860 1738 6 clka
rlabel metal2 532 1738 532 1738 6 clkb
rlabel metal3 2 1535 2 1535 6 reset
rlabel metal3 2 1205 2 1205 6 start
rlabel metal3 1765 1055 1765 1055 6 cordic_mode
rlabel metal3 1765 875 1765 875 6 in_port0[7]
rlabel metal3 1765 855 1765 855 6 in_port0[6]
rlabel metal3 1765 835 1765 835 6 in_port0[5]
rlabel metal3 1765 915 1765 915 6 in_port0[4]
rlabel metal3 1765 935 1765 935 6 in_port0[3]
rlabel metal3 1765 895 1765 895 6 in_port0[2]
rlabel metal3 1765 815 1765 815 6 in_port0[1]
rlabel metal2 972 1738 972 1738 6 in_port0[0]
rlabel metal3 2 1015 2 1015 6 in_port1[7]
rlabel metal3 2 925 2 925 6 in_port1[6]
rlabel metal3 2 995 2 995 6 in_port1[5]
rlabel metal3 2 815 2 815 6 in_port1[4]
rlabel metal3 2 615 2 615 6 in_port1[3]
rlabel metal3 2 525 2 525 6 in_port1[2]
rlabel metal3 2 325 2 325 6 in_port1[1]
rlabel metal3 2 305 2 305 6 in_port1[0]
rlabel metal3 1765 795 1765 795 6 out_port0[7]
rlabel metal3 1765 775 1765 775 6 out_port0[6]
rlabel metal3 1765 955 1765 955 6 out_port0[5]
rlabel metal3 1765 975 1765 975 6 out_port0[4]
rlabel metal3 1765 1015 1765 1015 6 out_port0[3]
rlabel metal3 1765 995 1765 995 6 out_port0[2]
rlabel metal3 1765 1035 1765 1035 6 out_port0[1]
rlabel metal2 988 1738 988 1738 6 out_port0[0]
rlabel metal2 732 1738 732 1738 6 out_port1[7]
rlabel metal3 2 905 2 905 6 out_port1[6]
rlabel metal3 2 1035 2 1035 6 out_port1[5]
rlabel metal3 2 795 2 795 6 out_port1[4]
rlabel metal3 2 675 2 675 6 out_port1[3]
rlabel metal3 2 475 2 475 6 out_port1[2]
rlabel metal3 2 275 2 275 6 out_port1[1]
rlabel metal3 2 225 2 225 6 out_port1[0]
rlabel metal2 420 1738 420 1738 6 done
rlabel metal1 38 367 38 367 6 gnd
rlabel metal1 14 67 14 67 6 vdd
<< end >>
