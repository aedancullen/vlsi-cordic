magic
tech scmos
timestamp 1683001453
<< metal1 >>
rect -1375 4088 -1314 4128
rect -1080 4097 -1019 4137
rect -778 4096 -717 4136
rect -482 4096 -421 4136
rect -170 4093 -109 4133
rect 121 4085 182 4125
rect 421 4086 470 4129
rect 715 4093 776 4133
rect 1023 4093 1084 4133
rect 1311 4085 1372 4125
rect 1621 4093 1682 4133
rect 1915 4085 1976 4125
rect -2232 3222 -2190 3282
rect -2230 2916 -2188 2976
rect 399 2740 498 3389
rect 918 3236 924 3304
rect 930 3236 936 3320
rect 942 3236 948 3288
rect 978 3107 984 3320
rect 990 3107 996 3263
rect 3981 3228 4021 3269
rect 1315 3207 1408 3215
rect 3992 2934 4032 2975
rect 894 2857 1020 2864
rect -2230 2629 -2188 2689
rect 3994 2641 4034 2682
rect -2232 2326 -2190 2386
rect -1491 2179 -945 2180
rect -1491 2177 -823 2179
rect -1491 2101 -839 2177
rect -824 2101 -823 2177
rect -1491 2099 -823 2101
rect -1491 2095 -945 2099
rect -2229 2021 -2189 2083
rect -1492 2060 -945 2095
rect -1492 2040 -1019 2060
rect -885 2051 -879 2056
rect -1492 2004 -1455 2040
rect -954 2012 -950 2016
rect -946 2012 -928 2016
rect -924 2012 -913 2016
rect -954 2011 -913 2012
rect -892 1925 -879 1926
rect -888 1921 -879 1925
rect -892 1815 -879 1816
rect -888 1811 -879 1815
rect 821 1791 894 1796
rect 900 1791 3293 1796
rect 821 1784 3293 1791
rect -2233 1716 -2191 1776
rect 821 1709 827 1784
rect 844 1709 3293 1784
rect 824 1708 3289 1709
rect -892 1695 -879 1696
rect -888 1691 -879 1695
rect -892 1495 -870 1496
rect -888 1491 -870 1495
rect -2232 1425 -2190 1485
rect -891 1295 -873 1296
rect -887 1291 -873 1295
rect -892 1245 -874 1246
rect -888 1241 -874 1245
rect -2229 1116 -2187 1176
rect -2229 825 -2187 885
rect -2226 523 -2184 583
rect -2235 -78 -2193 -18
rect -2228 -382 -2186 -322
rect -2229 -679 -2187 -619
rect -2225 -977 -2183 -917
rect -198 -1392 -97 1048
rect 22 -1378 111 -1374
rect 22 -1380 26 -1378
rect 111 -1390 115 -1378
rect -1077 -2134 -1029 -2092
rect -774 -2129 -726 -2087
rect -476 -2127 -428 -2085
rect 118 -2130 166 -2088
rect 429 -2130 477 -2088
rect 732 -2130 780 -2088
rect 1033 -2125 1081 -2083
rect 1331 -2127 1379 -2085
rect 1927 -2133 1975 -2091
rect 2231 -2136 2279 -2094
rect 2523 -2130 2571 -2088
<< m2contact >>
rect 3288 2910 3292 2915
rect 3285 2611 3289 2616
rect 3288 2311 3292 2315
rect -839 2101 -824 2177
rect -891 2051 -885 2056
rect 894 2051 900 2056
rect 894 2031 900 2037
rect -950 2012 -946 2016
rect -928 2012 -924 2016
rect 894 2011 900 2016
rect 894 1991 900 1996
rect 894 1971 900 1976
rect -892 1921 -888 1925
rect -892 1811 -888 1815
rect 894 1811 900 1816
rect 894 1791 900 1796
rect 827 1709 844 1784
rect -892 1691 -888 1695
rect -892 1491 -888 1495
rect -891 1291 -887 1295
rect -892 1241 -888 1245
rect -1493 -689 -1488 -685
rect -1491 -989 -1487 -985
rect -1494 -1289 -1488 -1285
rect -1389 -1393 -1385 -1387
rect -1089 -1392 -1085 -1386
rect -789 -1394 -785 -1388
rect 111 -1378 115 -1372
rect 22 -1386 26 -1380
rect 411 -1391 415 -1385
rect 711 -1394 715 -1388
rect 1011 -1393 1015 -1387
rect 1311 -1394 1315 -1388
rect 1910 -1395 1914 -1389
rect 2210 -1393 2214 -1387
<< metal2 >>
rect -1477 3378 -1471 3381
rect -1405 3378 -1399 3392
rect -1477 3372 -1399 3378
rect -1177 3368 -1171 3381
rect -1103 3368 -1097 3392
rect -1177 3362 -1097 3368
rect -877 3366 -871 3381
rect -805 3366 -799 3391
rect -877 3360 -799 3366
rect -577 3368 -571 3381
rect -506 3368 -500 3392
rect -577 3362 -500 3368
rect -277 3368 -271 3381
rect -204 3368 -198 3391
rect 23 3374 29 3381
rect 95 3374 101 3392
rect 23 3368 101 3374
rect 623 3369 629 3381
rect 694 3369 700 3392
rect -277 3362 -198 3368
rect 623 3363 700 3369
rect 923 3370 929 3381
rect 995 3370 1001 3392
rect 923 3364 1001 3370
rect 1223 3371 1229 3381
rect 1293 3371 1299 3391
rect 1223 3365 1299 3371
rect 1523 3366 1529 3381
rect 1597 3366 1603 3392
rect 1523 3360 1603 3366
rect 1823 3360 1829 3381
rect 1896 3360 1902 3392
rect 1823 3354 1902 3360
rect 930 3319 936 3320
rect 930 3313 931 3319
rect 935 3313 936 3319
rect 918 3303 924 3304
rect 918 3297 919 3303
rect 923 3297 924 3303
rect 918 3251 924 3297
rect 918 3238 919 3251
rect 923 3238 924 3251
rect 918 3236 924 3238
rect 930 3251 936 3313
rect 978 3319 984 3320
rect 978 3313 979 3319
rect 983 3313 984 3319
rect 930 3237 931 3251
rect 935 3237 936 3251
rect 930 3236 936 3237
rect 942 3287 948 3288
rect 942 3281 943 3287
rect 947 3281 948 3287
rect 942 3251 948 3281
rect 942 3237 943 3251
rect 947 3237 948 3251
rect 942 3236 948 3237
rect -1493 3193 -1467 3199
rect -1473 3129 -1467 3193
rect -1481 3123 -1467 3129
rect 978 3114 984 3313
rect 978 3108 979 3114
rect 983 3108 984 3114
rect 978 3107 984 3108
rect 990 3261 996 3263
rect 990 3252 991 3261
rect 995 3252 996 3261
rect 990 3114 996 3252
rect 1315 3214 1408 3215
rect 1315 3208 1316 3214
rect 1326 3208 1397 3214
rect 1407 3208 1408 3214
rect 1315 3207 1408 3208
rect 990 3108 991 3114
rect 995 3108 996 3114
rect 990 3107 996 3108
rect 3062 3149 3287 3152
rect -1481 3063 -1433 3066
rect -1481 3058 -1442 3063
rect -1437 3058 -1433 3063
rect -1481 3057 -1433 3058
rect -1445 3056 -1434 3057
rect -1492 2894 -1463 2900
rect -1469 2829 -1463 2894
rect 894 2863 1020 2864
rect 894 2858 895 2863
rect 899 2858 1009 2863
rect 1016 2858 1020 2863
rect 894 2857 1020 2858
rect -1482 2823 -1463 2829
rect 3062 2791 3065 3149
rect 3259 3123 3281 3129
rect 3259 2915 3265 3123
rect 3259 2910 3288 2915
rect 3259 2909 3292 2910
rect -442 2788 3065 2791
rect 3200 2849 3286 2852
rect -1481 2765 -1436 2766
rect -1481 2764 -1434 2765
rect -1481 2759 -1442 2764
rect -1436 2759 -1434 2764
rect -442 2761 -439 2788
rect 3200 2769 3203 2849
rect -150 2766 3203 2769
rect 3262 2823 3281 2829
rect -1481 2757 -1434 2759
rect -1445 2756 -1434 2757
rect -462 2752 -438 2761
rect -150 2755 -147 2766
rect 105 2756 3220 2761
rect -1493 2594 -1467 2600
rect -1473 2529 -1467 2594
rect 3215 2551 3220 2756
rect 3262 2616 3268 2823
rect 3262 2611 3285 2616
rect 3262 2610 3289 2611
rect 3215 2546 3286 2551
rect -1481 2523 -1467 2529
rect 3257 2523 3281 2529
rect -1481 2463 -1434 2466
rect -1481 2458 -1443 2463
rect -1437 2458 -1434 2463
rect -1481 2457 -1434 2458
rect -1445 2456 -1434 2457
rect 3257 2317 3263 2523
rect 3257 2315 3292 2317
rect 3257 2311 3288 2315
rect -1494 2296 -1462 2302
rect -1468 2229 -1462 2296
rect -1481 2223 -1462 2229
rect -1000 2051 -891 2056
rect 900 2051 972 2056
rect -1481 1871 -1468 1877
rect -1474 1807 -1468 1871
rect -1492 1801 -1468 1807
rect -1481 1642 -1435 1643
rect -1481 1640 -1434 1642
rect -1481 1635 -1438 1640
rect -1481 1634 -1434 1635
rect -1445 1633 -1434 1634
rect -1481 1565 -1435 1566
rect -1481 1563 -1434 1565
rect -1481 1558 -1442 1563
rect -1435 1558 -1434 1563
rect -1481 1557 -1434 1558
rect -1445 1556 -1434 1557
rect -1492 1393 -1465 1399
rect -1471 1329 -1465 1393
rect -1481 1323 -1465 1329
rect -1481 1263 -1434 1266
rect -1481 1258 -1443 1263
rect -1436 1258 -1434 1263
rect -1481 1257 -1434 1258
rect -1445 1256 -1434 1257
rect -1494 1093 -1464 1099
rect -1470 1029 -1464 1093
rect -1481 1023 -1464 1029
rect -1481 963 -1434 966
rect -1481 958 -1443 963
rect -1435 958 -1434 963
rect -1481 957 -1434 958
rect -1445 956 -1434 957
rect -1490 792 -1463 798
rect -1469 729 -1463 792
rect -1481 723 -1463 729
rect -1481 663 -1434 666
rect -1481 658 -1443 663
rect -1437 658 -1434 663
rect -1481 657 -1434 658
rect -1445 656 -1434 657
rect -1493 495 -1462 501
rect -1468 429 -1462 495
rect -1481 423 -1462 429
rect -1481 71 -1450 77
rect -1456 5 -1450 71
rect -1492 -1 -1450 5
rect -1000 -448 -994 2051
rect 900 2031 960 2037
rect 900 2011 948 2016
rect 900 1991 936 1996
rect 900 1971 924 1976
rect -1490 -454 -994 -448
rect -988 1921 -892 1926
rect -1481 -477 -1463 -471
rect -1469 -684 -1463 -477
rect -1493 -685 -1463 -684
rect -1488 -689 -1463 -685
rect -1493 -690 -1463 -689
rect -988 -749 -982 1921
rect -1488 -755 -982 -749
rect -976 1811 -892 1816
rect 900 1811 912 1816
rect -1481 -777 -1454 -771
rect -1460 -984 -1454 -777
rect -1492 -985 -1454 -984
rect -1492 -989 -1491 -985
rect -1487 -989 -1454 -985
rect -1492 -990 -1454 -989
rect -976 -1049 -970 1811
rect -1485 -1055 -970 -1049
rect -964 1691 -892 1696
rect -1481 -1077 -1465 -1071
rect -1471 -1284 -1465 -1077
rect -964 -1144 -958 1691
rect -1494 -1285 -1465 -1284
rect -1488 -1289 -1465 -1285
rect -1494 -1290 -1465 -1289
rect -1151 -1150 -958 -1144
rect -952 1491 -892 1496
rect -1390 -1371 -1171 -1365
rect -1390 -1387 -1384 -1371
rect -1177 -1381 -1171 -1371
rect -1390 -1393 -1389 -1387
rect -1385 -1393 -1384 -1387
rect -1151 -1389 -1145 -1150
rect -952 -1224 -946 1491
rect -940 1291 -891 1296
rect -940 -1191 -934 1291
rect -928 1241 -892 1246
rect -928 -1157 -922 1241
rect 894 -767 900 1791
rect 346 -773 900 -767
rect -928 -1163 47 -1157
rect -940 -1197 -555 -1191
rect -952 -1230 -844 -1224
rect -1091 -1374 -871 -1368
rect -1091 -1386 -1085 -1374
rect -877 -1382 -871 -1374
rect -850 -1384 -844 -1230
rect -791 -1377 -571 -1371
rect -1091 -1392 -1089 -1386
rect -791 -1388 -785 -1377
rect -577 -1381 -571 -1377
rect -561 -1382 -555 -1197
rect -561 -1388 -549 -1382
rect -791 -1394 -789 -1388
rect 41 -1391 47 -1163
rect 323 -1370 329 -1369
rect 109 -1372 329 -1370
rect 109 -1376 111 -1372
rect 110 -1378 111 -1376
rect 115 -1376 329 -1372
rect 115 -1378 116 -1376
rect 323 -1381 329 -1376
rect 346 -1390 352 -773
rect 906 -802 912 1811
rect 639 -808 912 -802
rect 410 -1374 629 -1368
rect 410 -1385 416 -1374
rect 623 -1381 629 -1374
rect 639 -1384 645 -808
rect 918 -848 924 1971
rect 930 -817 936 1991
rect 942 -787 948 2011
rect 954 -755 960 2031
rect 966 -716 972 2051
rect 966 -722 2450 -716
rect 954 -761 2148 -755
rect 942 -793 1848 -787
rect 930 -823 1263 -817
rect 918 -854 950 -848
rect 709 -1372 929 -1366
rect 410 -1391 411 -1385
rect 415 -1391 416 -1385
rect 410 -1392 416 -1391
rect 709 -1388 715 -1372
rect 923 -1384 929 -1372
rect 944 -1386 950 -854
rect 1011 -1376 1229 -1370
rect 709 -1394 711 -1388
rect 1011 -1387 1017 -1376
rect 1223 -1381 1229 -1376
rect 1015 -1393 1017 -1387
rect 1243 -1392 1249 -823
rect 1310 -1368 1829 -1362
rect 1310 -1388 1316 -1368
rect 1823 -1381 1829 -1368
rect 1310 -1394 1311 -1388
rect 1315 -1394 1316 -1388
rect 1842 -1389 1848 -793
rect 1909 -1374 2129 -1368
rect 1909 -1389 1915 -1374
rect 2123 -1382 2129 -1374
rect 2142 -1387 2148 -761
rect 2208 -1365 2429 -1359
rect 2208 -1387 2214 -1365
rect 2423 -1382 2429 -1365
rect 1909 -1395 1910 -1389
rect 1914 -1395 1915 -1389
rect 2208 -1393 2210 -1387
rect 2444 -1391 2450 -722
rect 1909 -1397 1915 -1395
<< m3contact >>
rect -1241 3379 -1234 3384
rect -940 3381 -936 3385
rect -1488 3359 -1484 3363
rect -640 3381 -636 3385
rect -339 3381 -335 3385
rect -39 3381 -35 3385
rect 261 3382 265 3387
rect 861 3381 865 3385
rect 1160 3381 1164 3385
rect 1459 3380 1463 3384
rect 1760 3381 1764 3385
rect 2057 3380 2061 3384
rect 931 3313 935 3319
rect 919 3297 923 3303
rect 919 3238 923 3251
rect 979 3313 983 3319
rect 931 3237 935 3251
rect 943 3281 947 3287
rect 943 3237 947 3251
rect 979 3108 983 3114
rect 991 3252 995 3261
rect 1316 3208 1326 3214
rect 1397 3208 1407 3214
rect 991 3108 995 3114
rect -1442 3058 -1437 3063
rect 895 2858 899 2863
rect 1009 2858 1016 2863
rect -1442 2759 -1436 2764
rect -350 2752 -346 2756
rect -22 2752 -18 2756
rect 90 2752 94 2756
rect -1443 2458 -1437 2463
rect -885 2052 -881 2056
rect 890 2052 894 2056
rect -1438 1635 -1434 1640
rect -1442 1558 -1435 1563
rect -1443 1258 -1436 1263
rect -1443 958 -1435 963
rect -1443 658 -1437 663
rect -1489 -164 -1482 -159
rect 890 2032 894 2036
rect -954 2012 -950 2016
rect -924 2012 -920 2016
rect 890 2012 894 2016
rect 890 1992 894 1996
rect 890 1972 894 1976
rect -888 1921 -884 1925
rect -888 1811 -884 1815
rect 890 1812 894 1816
rect 890 1792 894 1796
rect -888 1691 -884 1695
rect -888 1491 -884 1495
rect -887 1291 -883 1295
rect -888 1241 -884 1245
<< metal3 >>
rect 258 3387 267 3389
rect -942 3385 -933 3386
rect -1242 3384 -1233 3385
rect -1242 3379 -1241 3384
rect -1234 3379 -1233 3384
rect -1489 3363 -1324 3364
rect -1489 3359 -1488 3363
rect -1484 3359 -1324 3363
rect -1489 3358 -1324 3359
rect -1330 3195 -1324 3358
rect -1242 3225 -1233 3379
rect -942 3381 -940 3385
rect -936 3381 -933 3385
rect -942 3241 -933 3381
rect -642 3385 -633 3386
rect -642 3381 -640 3385
rect -636 3381 -633 3385
rect -642 3257 -633 3381
rect -342 3385 -333 3386
rect -342 3381 -339 3385
rect -335 3381 -333 3385
rect -342 3272 -333 3381
rect -42 3385 -33 3386
rect -42 3381 -39 3385
rect -35 3381 -33 3385
rect -42 3288 -33 3381
rect 258 3382 261 3387
rect 265 3382 267 3387
rect 258 3304 267 3382
rect 858 3385 867 3386
rect 858 3381 861 3385
rect 865 3381 867 3385
rect 858 3320 867 3381
rect 1158 3385 1167 3386
rect 1758 3385 1766 3386
rect 1158 3381 1160 3385
rect 1164 3381 1167 3385
rect 1158 3320 1167 3381
rect 1456 3384 1466 3385
rect 1456 3380 1459 3384
rect 1463 3380 1466 3384
rect 1456 3343 1466 3380
rect 1758 3381 1760 3385
rect 1764 3381 1766 3385
rect 858 3319 936 3320
rect 858 3313 931 3319
rect 935 3313 936 3319
rect 858 3312 936 3313
rect 978 3319 1167 3320
rect 978 3313 979 3319
rect 983 3313 1167 3319
rect 978 3312 1167 3313
rect 1365 3333 1468 3343
rect 258 3303 924 3304
rect 258 3297 919 3303
rect 923 3297 924 3303
rect 258 3296 924 3297
rect -42 3287 948 3288
rect -42 3281 943 3287
rect 947 3281 948 3287
rect -42 3280 948 3281
rect -343 3264 996 3272
rect 990 3261 996 3264
rect -642 3249 95 3257
rect 990 3252 991 3261
rect 995 3252 996 3261
rect -942 3233 -17 3241
rect -226 3232 -17 3233
rect -1242 3217 -345 3225
rect -1330 3185 -886 3195
rect -1445 3063 -898 3066
rect -1445 3058 -1442 3063
rect -1437 3058 -898 3063
rect -1445 3056 -898 3058
rect -1445 2764 -910 2766
rect -1445 2759 -1442 2764
rect -1436 2759 -910 2764
rect -1445 2756 -910 2759
rect -1445 2463 -934 2465
rect -1445 2458 -1443 2463
rect -1437 2458 -934 2463
rect -1445 2456 -934 2458
rect -955 2016 -949 2017
rect -1439 2012 -954 2016
rect -950 2012 -946 2016
rect -1439 2011 -946 2012
rect -1439 1640 -1433 2011
rect -940 1946 -934 2456
rect -916 2036 -910 2756
rect -904 2226 -898 3056
rect -892 2556 -886 3185
rect -351 2756 -345 3217
rect -22 2892 -17 3232
rect -351 2752 -350 2756
rect -346 2752 -345 2756
rect -351 2751 -345 2752
rect -23 2756 -17 2892
rect -23 2752 -22 2756
rect -18 2752 -17 2756
rect -23 2751 -17 2752
rect 89 2756 95 3249
rect 918 3251 924 3252
rect 918 3238 919 3251
rect 923 3238 924 3251
rect 89 2752 90 2756
rect 94 2752 95 2756
rect 89 2751 95 2752
rect 894 2863 900 2864
rect 894 2858 895 2863
rect 899 2858 900 2863
rect -892 2551 -866 2556
rect -904 2221 -866 2226
rect 894 2077 900 2858
rect 877 2071 900 2077
rect -886 2056 -880 2057
rect 889 2056 895 2057
rect -892 2052 -885 2056
rect -881 2052 -867 2056
rect -892 2051 -867 2052
rect 878 2052 890 2056
rect 894 2052 900 2056
rect 878 2051 900 2052
rect 877 2036 900 2037
rect -916 2031 -866 2036
rect 877 2032 890 2036
rect 894 2032 900 2036
rect 877 2031 900 2032
rect -925 2016 -919 2017
rect 889 2016 895 2017
rect -928 2012 -924 2016
rect -920 2012 -866 2016
rect -928 2011 -866 2012
rect 878 2012 890 2016
rect 894 2012 900 2016
rect 878 2011 900 2012
rect 889 1996 895 1997
rect 878 1992 890 1996
rect 894 1992 900 1996
rect 878 1991 900 1992
rect 889 1976 895 1977
rect 878 1972 890 1976
rect 894 1972 900 1976
rect 878 1971 900 1972
rect 918 1957 924 3238
rect 877 1951 924 1957
rect 930 3251 936 3252
rect 930 3237 931 3251
rect 935 3237 936 3251
rect -940 1941 -866 1946
rect 930 1937 936 3237
rect 877 1931 936 1937
rect 942 3251 948 3252
rect 990 3251 996 3252
rect 942 3237 943 3251
rect 947 3237 948 3251
rect -892 1925 -866 1926
rect -892 1921 -888 1925
rect -884 1921 -866 1925
rect -889 1920 -883 1921
rect 942 1917 948 3237
rect 878 1911 948 1917
rect 954 3214 1327 3215
rect 954 3208 1316 3214
rect 1326 3208 1327 3214
rect 954 3207 1327 3208
rect 954 1897 960 3207
rect 1365 3199 1375 3333
rect 1758 3215 1766 3381
rect 1396 3214 1766 3215
rect 1396 3208 1397 3214
rect 1407 3208 1766 3214
rect 1396 3207 1766 3208
rect 2055 3385 2060 3387
rect 2055 3384 2064 3385
rect 2055 3380 2057 3384
rect 2061 3380 2064 3384
rect 878 1891 960 1897
rect 966 3191 1375 3199
rect 966 1877 972 3191
rect 878 1871 972 1877
rect 978 3114 984 3119
rect 978 3108 979 3114
rect 983 3108 984 3114
rect 978 1857 984 3108
rect 882 1851 984 1857
rect 990 3114 996 3119
rect 990 3108 991 3114
rect 995 3108 996 3114
rect 990 1837 996 3108
rect 2055 3065 2064 3380
rect 1028 3056 2064 3065
rect 1028 2864 1034 3056
rect 1007 2863 1034 2864
rect 1007 2858 1009 2863
rect 1016 2858 1034 2863
rect 1007 2857 1034 2858
rect -1439 1635 -1438 1640
rect -1434 1635 -1433 1640
rect -1439 1633 -1433 1635
rect -1424 1831 -866 1836
rect 882 1831 996 1837
rect -1424 1565 -1418 1831
rect 889 1816 895 1817
rect -892 1815 -866 1816
rect -892 1811 -888 1815
rect -884 1811 -866 1815
rect 878 1812 890 1816
rect 894 1812 900 1816
rect 878 1811 900 1812
rect -889 1810 -883 1811
rect 889 1796 895 1797
rect 878 1792 890 1796
rect 894 1792 900 1796
rect 878 1791 900 1792
rect -892 1695 -866 1696
rect -892 1691 -888 1695
rect -884 1691 -866 1695
rect -889 1690 -883 1691
rect -1445 1563 -1418 1565
rect -1445 1558 -1442 1563
rect -1435 1558 -1418 1563
rect -1445 1556 -1418 1558
rect -1402 1631 -866 1636
rect -1402 1265 -1390 1631
rect -1445 1263 -1390 1265
rect -1445 1258 -1443 1263
rect -1436 1258 -1390 1263
rect -1445 1256 -1390 1258
rect -1370 1541 -866 1546
rect -1370 965 -1361 1541
rect -892 1495 -866 1496
rect -892 1491 -888 1495
rect -884 1491 -866 1495
rect -889 1490 -883 1491
rect -1445 963 -1361 965
rect -1445 958 -1443 963
rect -1435 958 -1361 963
rect -1445 956 -1361 958
rect -1334 1341 -866 1346
rect -1334 665 -1324 1341
rect -1445 663 -1324 665
rect -1445 658 -1443 663
rect -1437 658 -1324 663
rect -1445 656 -1324 658
rect -1299 1321 -866 1326
rect -1299 542 -1289 1321
rect -892 1295 -866 1296
rect -892 1291 -887 1295
rect -883 1291 -866 1295
rect -888 1290 -882 1291
rect -892 1245 -866 1246
rect -892 1241 -888 1245
rect -884 1241 -866 1245
rect -889 1240 -883 1241
rect -1299 530 -1233 542
rect -1242 -157 -1233 530
rect -1490 -159 -1233 -157
rect -1490 -164 -1489 -159
rect -1482 -164 -1233 -159
rect -1490 -166 -1233 -164
rect -1242 -171 -1233 -166
use PadFC  16_0
timestamp 1000338511
transform 1 0 -2500 0 1 3400
box 327 -3 1003 673
use PadBiDir  17_0
timestamp 1680926210
transform 1 0 -1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_1
timestamp 1680926210
transform 1 0 -1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_2
timestamp 1680926210
transform 1 0 -900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_3
timestamp 1680926210
transform 1 0 -600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_4
timestamp 1680926210
transform 1 0 -300 0 1 3400
box -36 -19 303 1000
use PadVdd  18_0
timestamp 1522810018
transform 1 0 300 0 1 3400
box -3 -12 303 1000
use PadBiDir  17_5
timestamp 1680926210
transform 1 0 0 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_6
timestamp 1680926210
transform 1 0 600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_7
timestamp 1680926210
transform 1 0 900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_8
timestamp 1680926210
transform 1 0 1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_0
timestamp 1680926210
transform 1 0 1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_1
timestamp 1680926210
transform 1 0 1800 0 1 3400
box -36 -19 303 1000
use PadVdd  PadVdd_0
timestamp 1522810018
transform 1 0 2400 0 1 3400
box -3 -12 303 1000
use PadBiDir  PadBiDir_2
timestamp 1680926210
transform 1 0 2100 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_3
timestamp 1680926210
transform 1 0 2700 0 1 3400
box -36 -19 303 1000
use PadFC  16_1
timestamp 1000338511
transform 0 1 3300 -1 0 4400
box 327 -3 1003 673
use PadBiDir  PadBiDir_4
timestamp 1680926210
transform 1 0 3000 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_9
timestamp 1680926210
transform 0 -1 -1500 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_10
timestamp 1680926210
transform 0 -1 -1500 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_17
timestamp 1680926210
transform 0 1 3300 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_18
timestamp 1680926210
transform 0 1 3300 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_11
timestamp 1680926210
transform 0 -1 -1500 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_12
timestamp 1680926210
transform 0 -1 -1500 1 0 2200
box -36 -19 303 1000
use PadGnd  19_0
timestamp 1522810115
transform 0 -1 -1500 -1 0 2200
box -3 -11 303 1000
use PadBiDir  17_13
timestamp 1680926210
transform 0 -1 -1500 -1 0 1900
box -36 -19 303 1000
use PadBiDir  PadBiDir_14
timestamp 1680926210
transform 0 -1 -1500 1 0 1300
box -36 -19 303 1000
use CORDIC_TOP  CORDIC_TOP_0
timestamp 1681696376
transform 1 0 -880 0 1 1019
box 0 13 1767 1740
use PadBiDir  17_19
timestamp 1680926210
transform 0 1 3300 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_20
timestamp 1680926210
transform 0 1 3300 1 0 2200
box -36 -19 303 1000
use PadBiDir  17_21
timestamp 1680926210
transform 0 1 3300 1 0 1900
box -36 -19 303 1000
use PadGnd  19_1
timestamp 1522810115
transform 0 1 3300 -1 0 1900
box -3 -11 303 1000
use PadBiDir  PadBiDir_19
timestamp 1680926210
transform 0 1 3300 1 0 1300
box -36 -19 303 1000
use PadBiDir  PadBiDir_13
timestamp 1680926210
transform 0 -1 -1500 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_12
timestamp 1680926210
transform 0 -1 -1500 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_11
timestamp 1680926210
transform 0 -1 -1500 1 0 400
box -36 -19 303 1000
use PadBiDir  PadBiDir_18
timestamp 1680926210
transform 0 1 3300 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_17
timestamp 1680926210
transform 0 1 3300 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_16
timestamp 1680926210
transform 0 1 3300 1 0 400
box -36 -19 303 1000
use PadGnd  PadGnd_0
timestamp 1522810115
transform 0 -1 -1500 -1 0 400
box -3 -11 303 1000
use PadBiDir  PadBiDir_15
timestamp 1680926210
transform 0 1 3300 1 0 100
box -36 -19 303 1000
use PadBiDir  PadBiDir_10
timestamp 1680926210
transform 0 -1 -1500 -1 0 100
box -36 -19 303 1000
use PadBiDir  17_14
timestamp 1680926210
transform 0 -1 -1500 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_15
timestamp 1680926210
transform 0 -1 -1500 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_16
timestamp 1680926210
transform 0 -1 -1500 1 0 -1100
box -36 -19 303 1000
use PadGnd  PadGnd_1
timestamp 1522810115
transform 0 1 3300 -1 0 100
box -3 -11 303 1000
use PadBiDir  17_22
timestamp 1680926210
transform 0 1 3300 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_23
timestamp 1680926210
transform 0 1 3300 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_24
timestamp 1680926210
transform 0 1 3300 1 0 -1100
box -36 -19 303 1000
use PadBiDir  17_25
timestamp 1680926210
transform 0 -1 -1500 1 0 -1400
box -36 -19 303 1000
use PadFC  16_2
timestamp 1000338511
transform 0 -1 -1500 1 0 -2400
box 327 -3 1003 673
use PadBiDir  17_26
timestamp 1680926210
transform 1 0 -1500 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_27
timestamp 1680926210
transform 1 0 -1200 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_28
timestamp 1680926210
transform 1 0 -900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_29
timestamp 1680926210
transform 1 0 -600 0 -1 -1400
box -36 -19 303 1000
use PadVdd  18_1
timestamp 1522810018
transform 1 0 -300 0 -1 -1400
box -3 -12 303 1000
use PadBiDir  17_30
timestamp 1680926210
transform 1 0 0 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_31
timestamp 1680926210
transform 1 0 300 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_32
timestamp 1680926210
transform 1 0 600 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_33
timestamp 1680926210
transform 1 0 900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_35
timestamp 1680926210
transform 1 0 1200 0 -1 -1400
box -36 -19 303 1000
use PadVdd  PadVdd_1
timestamp 1522810018
transform 1 0 1500 0 -1 -1400
box -3 -12 303 1000
use PadBiDir  PadBiDir_5
timestamp 1680926210
transform 1 0 1800 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_6
timestamp 1680926210
transform 1 0 2100 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_7
timestamp 1680926210
transform 1 0 2400 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_8
timestamp 1680926210
transform 1 0 2700 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_34
timestamp 1680926210
transform 0 1 3300 1 0 -1400
box -36 -19 303 1000
use PadFC  16_3
timestamp 1000338511
transform -1 0 4300 0 -1 -1400
box 327 -3 1003 673
use PadBiDir  PadBiDir_9
timestamp 1680926210
transform 1 0 3000 0 -1 -1400
box -36 -19 303 1000
<< labels >>
rlabel metal1 -1352 4113 -1352 4113 1 p_clkb
rlabel metal1 -1052 4111 -1052 4111 1 p_clka
rlabel metal1 -751 4115 -751 4115 1 p_in_port0_0
rlabel metal1 -455 4108 -455 4108 1 p_in_port0_1
rlabel metal1 -138 4113 -138 4113 1 p_in_port0_2
rlabel metal1 149 4102 149 4102 1 p_in_port0_3
rlabel metal1 739 4111 739 4111 1 p_in_port0_4
rlabel metal1 1046 4120 1046 4120 1 p_in_port0_5
rlabel metal1 1334 4104 1334 4104 1 p_in_port0_6
rlabel metal1 1652 4117 1652 4117 1 p_in_port0_7
rlabel metal1 1940 4100 1940 4100 1 p_cordic_mode
rlabel metal1 -2208 2655 -2208 2655 1 p_in_port1_7
rlabel metal1 -2210 2357 -2210 2357 1 p_in_port1_6
rlabel metal1 -2217 1746 -2217 1746 1 p_in_port1_5
rlabel metal1 -2215 1447 -2215 1447 1 p_in_port1_4
rlabel metal1 -2208 1156 -2208 1156 1 p_in_port1_3
rlabel metal1 -2204 843 -2204 843 1 p_in_port1_2
rlabel metal1 -2208 550 -2208 550 1 p_in_port1_1
rlabel metal1 -2217 -41 -2217 -41 1 p_in_port1_0
rlabel metal1 -2204 -354 -2204 -354 1 p_out_port1_5
rlabel metal1 -2208 -656 -2208 -656 1 p_out_port1_6
rlabel metal1 -2204 -945 -2204 -945 1 p_out_port1_4
rlabel metal1 -1047 -2110 -1047 -2110 1 p_out_port1_3
rlabel metal1 -750 -2106 -750 -2106 1 p_out_port1_2
rlabel metal1 -455 -2108 -455 -2108 1 p_out_port1_1
rlabel metal1 138 -2103 138 -2103 1 p_out_port1_0
rlabel metal1 456 -2106 456 -2106 1 p_out_port0_6
rlabel metal1 751 -2115 751 -2115 1 p_out_port0_7
rlabel metal1 1055 -2106 1055 -2106 1 p_out_port0_5
rlabel metal1 1364 -2103 1364 -2103 1 p_out_port0_4
rlabel metal1 1939 -2108 1939 -2108 1 p_out_port0_2
rlabel metal1 2250 -2110 2250 -2110 1 p_out_port0_3
rlabel metal1 2541 -2106 2541 -2106 1 p_out_port0_1
rlabel metal1 4002 3255 4002 3255 1 p_done
rlabel metal1 4007 2957 4007 2957 1 p_out_port1_7
rlabel metal1 4016 2663 4016 2663 1 p_out_port0_0
rlabel metal1 -2210 3254 -2210 3254 1 p_reset
rlabel metal1 -2213 2945 -2213 2945 1 p_start
rlabel metal2 909 1974 909 1974 1 out_port0_5
rlabel metal1 446 4106 446 4106 1 Vdd
rlabel metal1 -2210 2051 -2210 2051 1 GND
rlabel metal3 903 1833 903 1833 1 in_port0_1
rlabel metal3 903 1854 903 1854 1 in_port0_5
rlabel metal3 902 1873 902 1873 1 in_port0_6
rlabel metal3 900 1894 900 1894 1 in_port0_7
rlabel metal3 899 1912 899 1912 1 in_port0_2
rlabel metal3 899 1933 899 1933 1 in_port0_4
rlabel metal3 899 1954 899 1954 1 in_port0_3
rlabel metal3 896 2074 896 2074 1 cordic_mode
rlabel m3contact -348 2753 -348 2753 1 clkb
rlabel m3contact 92 2754 92 2754 1 in_port0_0
rlabel m3contact -20 2753 -20 2753 1 clka
rlabel metal3 -873 2554 -873 2554 1 reset
rlabel metal3 -872 2223 -872 2223 1 start
rlabel metal3 -870 2033 -870 2033 1 in_port1_7
rlabel metal3 -870 2014 -870 2014 1 in_port1_5
rlabel metal3 -870 1943 -870 1943 1 in_port1_6
rlabel metal3 -870 1833 -870 1833 1 in_port1_4
rlabel metal3 -869 1632 -869 1632 1 in_port1_3
rlabel metal3 -869 1543 -869 1543 1 in_port1_2
rlabel metal3 -869 1343 -869 1343 1 in_port1_1
rlabel metal3 -868 1324 -868 1324 1 in_port1_0
<< end >>
