magic
tech scmos
timestamp 1683038052
<< nwell >>
rect -9 48 26 105
<< ntransistor >>
rect 7 6 9 26
<< ptransistor >>
rect 7 54 9 94
<< ndiffusion >>
rect 2 6 7 26
rect 9 6 14 26
<< pdiffusion >>
rect 2 54 7 94
rect 9 54 14 94
<< psubstratepdiff >>
rect -2 -2 2 2
<< nsubstratendiff >>
rect -2 98 2 102
<< polysilicon >>
rect 7 94 9 96
rect 7 33 9 54
rect 2 29 9 33
rect 7 26 9 29
rect 7 4 9 6
<< genericcontact >>
rect -1 99 1 101
rect 3 90 5 92
rect 11 90 13 92
rect 3 85 5 87
rect 11 85 13 87
rect 3 80 5 82
rect 11 80 13 82
rect 3 75 5 77
rect 11 75 13 77
rect 3 70 5 72
rect 11 70 13 72
rect 3 65 5 67
rect 11 65 13 67
rect 3 60 5 62
rect 11 60 13 62
rect 3 55 5 57
rect 11 55 13 57
rect 3 30 5 32
rect 3 22 5 24
rect 11 22 13 24
rect 3 17 5 19
rect 11 17 13 19
rect 3 12 5 14
rect 11 12 13 14
rect 3 7 5 9
rect 11 7 13 9
rect -1 -1 1 1
<< metal1 >>
rect -2 97 18 103
rect 2 54 6 97
rect 2 29 6 37
rect 2 3 6 26
rect 10 6 14 94
rect -2 -3 18 3
<< m1p >>
rect 10 43 14 47
rect 2 33 6 37
<< labels >>
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 12 45 12 45 6 Y
rlabel metal1 4 35 4 35 6 A
<< end >>
