magic
tech scmos
timestamp 1683038052
<< nwell >>
rect 20 740 280 1000
rect 17 429 283 653
rect -3 249 303 330
rect -3 11 11 249
rect 289 11 303 249
rect -3 -3 303 11
<< ptransistor >>
rect 38 626 138 629
rect 38 582 138 585
rect 38 562 138 565
rect 38 518 138 521
rect 38 497 138 500
rect 38 453 138 456
rect 162 626 262 629
rect 162 582 262 585
rect 162 562 262 565
rect 162 518 262 521
rect 162 497 262 500
rect 162 453 262 456
<< pdiffusion >>
rect 38 629 138 638
rect 38 585 138 626
rect 38 565 138 582
rect 38 521 138 562
rect 38 500 138 518
rect 38 456 138 497
rect 38 444 138 453
rect 162 629 262 638
rect 162 585 262 626
rect 162 565 262 582
rect 162 521 262 562
rect 162 500 262 518
rect 162 456 262 497
rect 162 444 262 453
<< psubstratepdiff >>
rect 0 659 300 670
rect 0 423 11 659
rect 289 423 300 659
rect 0 343 300 423
rect 14 14 286 246
<< nsubstratendiff >>
rect 20 640 280 650
rect 20 442 30 640
rect 36 638 138 640
rect 38 442 138 444
rect 142 442 158 640
rect 162 638 264 640
rect 162 442 262 444
rect 270 442 280 640
rect 20 432 280 442
rect 0 252 300 327
rect 0 8 8 252
rect 292 8 300 252
rect 0 0 300 8
<< polysilicon >>
rect 2 715 17 718
rect 20 715 35 718
rect 8 703 11 715
rect 20 712 23 715
rect 32 712 35 715
rect 20 709 35 712
rect 20 703 23 709
rect 32 703 35 709
rect 38 715 41 718
rect 38 712 47 715
rect 38 703 41 712
rect 44 709 47 712
rect 50 709 53 718
rect 44 706 53 709
rect 50 703 53 706
rect 56 715 59 718
rect 56 712 65 715
rect 56 703 59 712
rect 62 709 65 712
rect 68 709 71 718
rect 62 706 71 709
rect 68 703 71 706
rect 74 715 89 718
rect 92 715 107 718
rect 74 712 77 715
rect 92 712 95 715
rect 104 712 107 715
rect 74 709 89 712
rect 92 709 107 712
rect 74 706 77 709
rect 74 703 89 706
rect 92 703 95 709
rect 101 703 104 709
rect 194 707 209 710
rect 194 695 197 707
rect 200 701 203 707
rect 206 695 209 707
rect 212 707 227 710
rect 212 698 215 707
rect 224 698 227 707
rect 230 707 245 710
rect 248 707 263 710
rect 266 707 281 710
rect 230 704 233 707
rect 230 701 245 704
rect 242 698 245 701
rect 254 698 257 707
rect 266 704 269 707
rect 266 701 281 704
rect 278 698 281 701
rect 212 695 227 698
rect 230 695 245 698
rect 248 695 263 698
rect 266 695 281 698
rect 42 689 57 692
rect 60 689 75 692
rect 78 689 93 692
rect 42 680 45 689
rect 60 686 63 689
rect 78 686 81 689
rect 60 683 75 686
rect 78 683 93 686
rect 60 680 63 683
rect 90 680 93 683
rect 42 677 57 680
rect 60 677 75 680
rect 78 677 93 680
rect 31 626 38 629
rect 138 626 140 629
rect 31 585 37 626
rect 31 582 38 585
rect 138 582 140 585
rect 31 565 37 582
rect 31 562 38 565
rect 138 562 140 565
rect 31 521 37 562
rect 31 518 38 521
rect 138 518 140 521
rect 31 500 37 518
rect 31 497 38 500
rect 138 497 140 500
rect 31 456 37 497
rect 31 453 38 456
rect 138 453 140 456
rect 160 626 162 629
rect 262 626 269 629
rect 263 585 269 626
rect 160 582 162 585
rect 262 582 269 585
rect 263 565 269 582
rect 160 562 162 565
rect 262 562 269 565
rect 263 521 269 562
rect 160 518 162 521
rect 262 518 269 521
rect 263 500 269 518
rect 160 497 162 500
rect 262 497 269 500
rect 263 456 269 497
rect 160 453 162 456
rect 262 453 269 456
<< genericcontact >>
rect 2 666 4 668
rect 7 666 9 668
rect 12 666 14 668
rect 17 666 19 668
rect 22 666 24 668
rect 27 666 29 668
rect 32 666 34 668
rect 37 666 39 668
rect 42 666 44 668
rect 47 666 49 668
rect 52 666 54 668
rect 57 666 59 668
rect 62 666 64 668
rect 67 666 69 668
rect 72 666 74 668
rect 77 666 79 668
rect 82 666 84 668
rect 87 666 89 668
rect 92 666 94 668
rect 97 666 99 668
rect 102 666 104 668
rect 107 666 109 668
rect 112 666 114 668
rect 117 666 119 668
rect 122 666 124 668
rect 127 666 129 668
rect 171 666 173 668
rect 176 666 178 668
rect 181 666 183 668
rect 186 666 188 668
rect 191 666 193 668
rect 196 666 198 668
rect 201 666 203 668
rect 206 666 208 668
rect 211 666 213 668
rect 216 666 218 668
rect 221 666 223 668
rect 226 666 228 668
rect 231 666 233 668
rect 236 666 238 668
rect 241 666 243 668
rect 246 666 248 668
rect 251 666 253 668
rect 256 666 258 668
rect 261 666 263 668
rect 266 666 268 668
rect 271 666 273 668
rect 276 666 278 668
rect 281 666 283 668
rect 286 666 288 668
rect 291 666 293 668
rect 296 666 298 668
rect 2 661 4 663
rect 7 661 9 663
rect 12 661 14 663
rect 17 661 19 663
rect 22 661 24 663
rect 27 661 29 663
rect 32 661 34 663
rect 37 661 39 663
rect 42 661 44 663
rect 47 661 49 663
rect 52 661 54 663
rect 57 661 59 663
rect 62 661 64 663
rect 67 661 69 663
rect 72 661 74 663
rect 77 661 79 663
rect 82 661 84 663
rect 87 661 89 663
rect 92 661 94 663
rect 97 661 99 663
rect 102 661 104 663
rect 107 661 109 663
rect 112 661 114 663
rect 117 661 119 663
rect 122 661 124 663
rect 127 661 129 663
rect 171 661 173 663
rect 176 661 178 663
rect 181 661 183 663
rect 186 661 188 663
rect 191 661 193 663
rect 196 661 198 663
rect 201 661 203 663
rect 206 661 208 663
rect 211 661 213 663
rect 216 661 218 663
rect 221 661 223 663
rect 226 661 228 663
rect 231 661 233 663
rect 236 661 238 663
rect 241 661 243 663
rect 246 661 248 663
rect 251 661 253 663
rect 256 661 258 663
rect 261 661 263 663
rect 266 661 268 663
rect 271 661 273 663
rect 276 661 278 663
rect 281 661 283 663
rect 286 661 288 663
rect 291 661 293 663
rect 296 661 298 663
rect 2 655 4 657
rect 7 655 9 657
rect 291 655 293 657
rect 296 655 298 657
rect 2 650 4 652
rect 7 650 9 652
rect 291 650 293 652
rect 296 650 298 652
rect 2 645 4 647
rect 7 645 9 647
rect 27 646 29 648
rect 271 646 273 648
rect 37 644 39 646
rect 42 644 44 646
rect 47 644 49 646
rect 52 644 54 646
rect 57 644 59 646
rect 62 644 64 646
rect 67 644 69 646
rect 72 644 74 646
rect 77 644 79 646
rect 82 644 84 646
rect 87 644 89 646
rect 92 644 94 646
rect 97 644 99 646
rect 102 644 104 646
rect 107 644 109 646
rect 112 644 114 646
rect 117 644 119 646
rect 181 644 183 646
rect 186 644 188 646
rect 191 644 193 646
rect 196 644 198 646
rect 201 644 203 646
rect 206 644 208 646
rect 211 644 213 646
rect 216 644 218 646
rect 221 644 223 646
rect 226 644 228 646
rect 231 644 233 646
rect 236 644 238 646
rect 241 644 243 646
rect 246 644 248 646
rect 251 644 253 646
rect 256 644 258 646
rect 261 644 263 646
rect 291 645 293 647
rect 296 645 298 647
rect 2 640 4 642
rect 7 640 9 642
rect 27 641 29 643
rect 271 641 273 643
rect 291 640 293 642
rect 296 640 298 642
rect 2 635 4 637
rect 7 635 9 637
rect 27 636 29 638
rect 271 636 273 638
rect 291 635 293 637
rect 296 635 298 637
rect 42 633 44 635
rect 47 633 49 635
rect 52 633 54 635
rect 57 633 59 635
rect 62 633 64 635
rect 67 633 69 635
rect 72 633 74 635
rect 77 633 79 635
rect 82 633 84 635
rect 87 633 89 635
rect 92 633 94 635
rect 97 633 99 635
rect 102 633 104 635
rect 107 633 109 635
rect 112 633 114 635
rect 117 633 119 635
rect 181 633 183 635
rect 186 633 188 635
rect 191 633 193 635
rect 196 633 198 635
rect 201 633 203 635
rect 206 633 208 635
rect 211 633 213 635
rect 216 633 218 635
rect 221 633 223 635
rect 226 633 228 635
rect 231 633 233 635
rect 236 633 238 635
rect 241 633 243 635
rect 246 633 248 635
rect 251 633 253 635
rect 256 633 258 635
rect 2 630 4 632
rect 7 630 9 632
rect 27 631 29 633
rect 271 631 273 633
rect 291 630 293 632
rect 296 630 298 632
rect 2 625 4 627
rect 7 625 9 627
rect 27 626 29 628
rect 271 626 273 628
rect 291 625 293 627
rect 296 625 298 627
rect 33 623 35 625
rect 265 623 267 625
rect 2 620 4 622
rect 7 620 9 622
rect 27 621 29 623
rect 271 621 273 623
rect 291 620 293 622
rect 296 620 298 622
rect 33 618 35 620
rect 265 618 267 620
rect 2 615 4 617
rect 7 615 9 617
rect 27 616 29 618
rect 271 616 273 618
rect 291 615 293 617
rect 296 615 298 617
rect 33 613 35 615
rect 2 610 4 612
rect 7 610 9 612
rect 27 611 29 613
rect 144 612 146 614
rect 149 612 151 614
rect 154 612 156 614
rect 265 613 267 615
rect 271 611 273 613
rect 291 610 293 612
rect 296 610 298 612
rect 33 608 35 610
rect 2 605 4 607
rect 7 605 9 607
rect 27 606 29 608
rect 57 607 59 609
rect 62 607 64 609
rect 67 607 69 609
rect 72 607 74 609
rect 77 607 79 609
rect 82 607 84 609
rect 87 607 89 609
rect 92 607 94 609
rect 97 607 99 609
rect 102 607 104 609
rect 107 607 109 609
rect 112 607 114 609
rect 117 607 119 609
rect 181 607 183 609
rect 186 607 188 609
rect 191 607 193 609
rect 196 607 198 609
rect 201 607 203 609
rect 206 607 208 609
rect 211 607 213 609
rect 216 607 218 609
rect 221 607 223 609
rect 226 607 228 609
rect 231 607 233 609
rect 236 607 238 609
rect 241 607 243 609
rect 265 608 267 610
rect 271 606 273 608
rect 291 605 293 607
rect 296 605 298 607
rect 33 603 35 605
rect 2 600 4 602
rect 7 600 9 602
rect 27 601 29 603
rect 57 602 59 604
rect 62 602 64 604
rect 67 602 69 604
rect 72 602 74 604
rect 77 602 79 604
rect 82 602 84 604
rect 87 602 89 604
rect 92 602 94 604
rect 97 602 99 604
rect 102 602 104 604
rect 107 602 109 604
rect 112 602 114 604
rect 117 602 119 604
rect 144 602 146 604
rect 149 602 151 604
rect 154 602 156 604
rect 181 602 183 604
rect 186 602 188 604
rect 191 602 193 604
rect 196 602 198 604
rect 201 602 203 604
rect 206 602 208 604
rect 211 602 213 604
rect 216 602 218 604
rect 221 602 223 604
rect 226 602 228 604
rect 231 602 233 604
rect 236 602 238 604
rect 241 602 243 604
rect 265 603 267 605
rect 271 601 273 603
rect 291 600 293 602
rect 296 600 298 602
rect 33 598 35 600
rect 265 598 267 600
rect 2 595 4 597
rect 7 595 9 597
rect 27 596 29 598
rect 271 596 273 598
rect 291 595 293 597
rect 296 595 298 597
rect 33 593 35 595
rect 2 590 4 592
rect 7 590 9 592
rect 27 591 29 593
rect 144 592 146 594
rect 149 592 151 594
rect 154 592 156 594
rect 265 593 267 595
rect 271 591 273 593
rect 291 590 293 592
rect 296 590 298 592
rect 33 588 35 590
rect 265 588 267 590
rect 2 585 4 587
rect 7 585 9 587
rect 27 586 29 588
rect 271 586 273 588
rect 291 585 293 587
rect 296 585 298 587
rect 33 583 35 585
rect 265 583 267 585
rect 2 580 4 582
rect 7 580 9 582
rect 27 581 29 583
rect 271 581 273 583
rect 291 580 293 582
rect 296 580 298 582
rect 33 578 35 580
rect 265 578 267 580
rect 2 575 4 577
rect 7 575 9 577
rect 27 576 29 578
rect 42 575 44 577
rect 47 575 49 577
rect 52 575 54 577
rect 57 575 59 577
rect 62 575 64 577
rect 67 575 69 577
rect 72 575 74 577
rect 77 575 79 577
rect 82 575 84 577
rect 87 575 89 577
rect 92 575 94 577
rect 97 575 99 577
rect 102 575 104 577
rect 107 575 109 577
rect 112 575 114 577
rect 117 575 119 577
rect 181 575 183 577
rect 186 575 188 577
rect 191 575 193 577
rect 196 575 198 577
rect 201 575 203 577
rect 206 575 208 577
rect 211 575 213 577
rect 216 575 218 577
rect 221 575 223 577
rect 226 575 228 577
rect 231 575 233 577
rect 236 575 238 577
rect 241 575 243 577
rect 246 575 248 577
rect 251 575 253 577
rect 256 575 258 577
rect 271 576 273 578
rect 291 575 293 577
rect 296 575 298 577
rect 33 573 35 575
rect 265 573 267 575
rect 2 570 4 572
rect 7 570 9 572
rect 27 571 29 573
rect 42 570 44 572
rect 47 570 49 572
rect 52 570 54 572
rect 57 570 59 572
rect 62 570 64 572
rect 67 570 69 572
rect 72 570 74 572
rect 77 570 79 572
rect 82 570 84 572
rect 87 570 89 572
rect 92 570 94 572
rect 97 570 99 572
rect 102 570 104 572
rect 107 570 109 572
rect 112 570 114 572
rect 117 570 119 572
rect 181 570 183 572
rect 186 570 188 572
rect 191 570 193 572
rect 196 570 198 572
rect 201 570 203 572
rect 206 570 208 572
rect 211 570 213 572
rect 216 570 218 572
rect 221 570 223 572
rect 226 570 228 572
rect 231 570 233 572
rect 236 570 238 572
rect 241 570 243 572
rect 246 570 248 572
rect 251 570 253 572
rect 256 570 258 572
rect 271 571 273 573
rect 291 570 293 572
rect 296 570 298 572
rect 33 568 35 570
rect 265 568 267 570
rect 2 565 4 567
rect 7 565 9 567
rect 27 566 29 568
rect 271 566 273 568
rect 291 565 293 567
rect 296 565 298 567
rect 33 563 35 565
rect 265 563 267 565
rect 2 560 4 562
rect 7 560 9 562
rect 27 561 29 563
rect 271 561 273 563
rect 291 560 293 562
rect 296 560 298 562
rect 33 558 35 560
rect 265 558 267 560
rect 2 555 4 557
rect 7 555 9 557
rect 27 556 29 558
rect 271 556 273 558
rect 291 555 293 557
rect 296 555 298 557
rect 33 553 35 555
rect 265 553 267 555
rect 2 550 4 552
rect 7 550 9 552
rect 27 551 29 553
rect 271 551 273 553
rect 291 550 293 552
rect 296 550 298 552
rect 33 548 35 550
rect 144 548 146 550
rect 149 548 151 550
rect 154 548 156 550
rect 265 548 267 550
rect 2 545 4 547
rect 7 545 9 547
rect 27 546 29 548
rect 271 546 273 548
rect 291 545 293 547
rect 296 545 298 547
rect 33 543 35 545
rect 57 543 59 545
rect 62 543 64 545
rect 67 543 69 545
rect 72 543 74 545
rect 77 543 79 545
rect 82 543 84 545
rect 87 543 89 545
rect 92 543 94 545
rect 97 543 99 545
rect 102 543 104 545
rect 107 543 109 545
rect 112 543 114 545
rect 117 543 119 545
rect 181 543 183 545
rect 186 543 188 545
rect 191 543 193 545
rect 196 543 198 545
rect 201 543 203 545
rect 206 543 208 545
rect 211 543 213 545
rect 216 543 218 545
rect 221 543 223 545
rect 226 543 228 545
rect 231 543 233 545
rect 236 543 238 545
rect 241 543 243 545
rect 265 543 267 545
rect 2 540 4 542
rect 7 540 9 542
rect 27 541 29 543
rect 271 541 273 543
rect 291 540 293 542
rect 296 540 298 542
rect 33 538 35 540
rect 57 538 59 540
rect 62 538 64 540
rect 67 538 69 540
rect 72 538 74 540
rect 77 538 79 540
rect 82 538 84 540
rect 87 538 89 540
rect 92 538 94 540
rect 97 538 99 540
rect 102 538 104 540
rect 107 538 109 540
rect 112 538 114 540
rect 117 538 119 540
rect 144 538 146 540
rect 149 538 151 540
rect 154 538 156 540
rect 181 538 183 540
rect 186 538 188 540
rect 191 538 193 540
rect 196 538 198 540
rect 201 538 203 540
rect 206 538 208 540
rect 211 538 213 540
rect 216 538 218 540
rect 221 538 223 540
rect 226 538 228 540
rect 231 538 233 540
rect 236 538 238 540
rect 241 538 243 540
rect 265 538 267 540
rect 2 535 4 537
rect 7 535 9 537
rect 27 536 29 538
rect 271 536 273 538
rect 291 535 293 537
rect 296 535 298 537
rect 33 533 35 535
rect 265 533 267 535
rect 2 530 4 532
rect 7 530 9 532
rect 27 531 29 533
rect 271 531 273 533
rect 291 530 293 532
rect 296 530 298 532
rect 33 528 35 530
rect 144 528 146 530
rect 149 528 151 530
rect 154 528 156 530
rect 265 528 267 530
rect 2 525 4 527
rect 7 525 9 527
rect 27 526 29 528
rect 271 526 273 528
rect 291 525 293 527
rect 296 525 298 527
rect 33 523 35 525
rect 265 523 267 525
rect 2 520 4 522
rect 7 520 9 522
rect 27 521 29 523
rect 271 521 273 523
rect 291 520 293 522
rect 296 520 298 522
rect 33 518 35 520
rect 265 518 267 520
rect 2 515 4 517
rect 7 515 9 517
rect 27 516 29 518
rect 271 516 273 518
rect 291 515 293 517
rect 296 515 298 517
rect 33 513 35 515
rect 265 513 267 515
rect 2 510 4 512
rect 7 510 9 512
rect 27 511 29 513
rect 42 511 44 513
rect 47 511 49 513
rect 52 511 54 513
rect 57 511 59 513
rect 62 511 64 513
rect 67 511 69 513
rect 72 511 74 513
rect 77 511 79 513
rect 82 511 84 513
rect 87 511 89 513
rect 92 511 94 513
rect 97 511 99 513
rect 102 511 104 513
rect 107 511 109 513
rect 112 511 114 513
rect 117 511 119 513
rect 181 511 183 513
rect 186 511 188 513
rect 191 511 193 513
rect 196 511 198 513
rect 201 511 203 513
rect 206 511 208 513
rect 211 511 213 513
rect 216 511 218 513
rect 221 511 223 513
rect 226 511 228 513
rect 231 511 233 513
rect 236 511 238 513
rect 241 511 243 513
rect 246 511 248 513
rect 251 511 253 513
rect 256 511 258 513
rect 271 511 273 513
rect 291 510 293 512
rect 296 510 298 512
rect 33 508 35 510
rect 265 508 267 510
rect 2 505 4 507
rect 7 505 9 507
rect 27 506 29 508
rect 42 505 44 507
rect 47 505 49 507
rect 52 505 54 507
rect 57 505 59 507
rect 62 505 64 507
rect 67 505 69 507
rect 72 505 74 507
rect 77 505 79 507
rect 82 505 84 507
rect 87 505 89 507
rect 92 505 94 507
rect 97 505 99 507
rect 102 505 104 507
rect 107 505 109 507
rect 112 505 114 507
rect 117 505 119 507
rect 181 505 183 507
rect 186 505 188 507
rect 191 505 193 507
rect 196 505 198 507
rect 201 505 203 507
rect 206 505 208 507
rect 211 505 213 507
rect 216 505 218 507
rect 221 505 223 507
rect 226 505 228 507
rect 231 505 233 507
rect 236 505 238 507
rect 241 505 243 507
rect 246 505 248 507
rect 251 505 253 507
rect 256 505 258 507
rect 271 506 273 508
rect 291 505 293 507
rect 296 505 298 507
rect 33 503 35 505
rect 265 503 267 505
rect 2 500 4 502
rect 7 500 9 502
rect 27 501 29 503
rect 271 501 273 503
rect 291 500 293 502
rect 296 500 298 502
rect 33 498 35 500
rect 265 498 267 500
rect 2 495 4 497
rect 7 495 9 497
rect 27 496 29 498
rect 271 496 273 498
rect 291 495 293 497
rect 296 495 298 497
rect 33 493 35 495
rect 265 493 267 495
rect 2 490 4 492
rect 7 490 9 492
rect 27 491 29 493
rect 271 491 273 493
rect 291 490 293 492
rect 296 490 298 492
rect 33 488 35 490
rect 265 488 267 490
rect 2 485 4 487
rect 7 485 9 487
rect 27 486 29 488
rect 271 486 273 488
rect 291 485 293 487
rect 296 485 298 487
rect 33 483 35 485
rect 144 483 146 485
rect 149 483 151 485
rect 154 483 156 485
rect 265 483 267 485
rect 2 480 4 482
rect 7 480 9 482
rect 27 481 29 483
rect 271 481 273 483
rect 291 480 293 482
rect 296 480 298 482
rect 33 478 35 480
rect 57 478 59 480
rect 62 478 64 480
rect 67 478 69 480
rect 72 478 74 480
rect 77 478 79 480
rect 82 478 84 480
rect 87 478 89 480
rect 92 478 94 480
rect 97 478 99 480
rect 102 478 104 480
rect 107 478 109 480
rect 112 478 114 480
rect 117 478 119 480
rect 181 478 183 480
rect 186 478 188 480
rect 191 478 193 480
rect 196 478 198 480
rect 201 478 203 480
rect 206 478 208 480
rect 211 478 213 480
rect 216 478 218 480
rect 221 478 223 480
rect 226 478 228 480
rect 231 478 233 480
rect 236 478 238 480
rect 241 478 243 480
rect 265 478 267 480
rect 2 475 4 477
rect 7 475 9 477
rect 27 476 29 478
rect 271 476 273 478
rect 291 475 293 477
rect 296 475 298 477
rect 33 473 35 475
rect 57 473 59 475
rect 62 473 64 475
rect 67 473 69 475
rect 72 473 74 475
rect 77 473 79 475
rect 82 473 84 475
rect 87 473 89 475
rect 92 473 94 475
rect 97 473 99 475
rect 102 473 104 475
rect 107 473 109 475
rect 112 473 114 475
rect 117 473 119 475
rect 144 473 146 475
rect 149 473 151 475
rect 154 473 156 475
rect 181 473 183 475
rect 186 473 188 475
rect 191 473 193 475
rect 196 473 198 475
rect 201 473 203 475
rect 206 473 208 475
rect 211 473 213 475
rect 216 473 218 475
rect 221 473 223 475
rect 226 473 228 475
rect 231 473 233 475
rect 236 473 238 475
rect 241 473 243 475
rect 265 473 267 475
rect 2 470 4 472
rect 7 470 9 472
rect 27 471 29 473
rect 271 471 273 473
rect 291 470 293 472
rect 296 470 298 472
rect 33 468 35 470
rect 265 468 267 470
rect 2 465 4 467
rect 7 465 9 467
rect 27 466 29 468
rect 271 466 273 468
rect 291 465 293 467
rect 296 465 298 467
rect 33 463 35 465
rect 144 463 146 465
rect 149 463 151 465
rect 154 463 156 465
rect 265 463 267 465
rect 2 460 4 462
rect 7 460 9 462
rect 27 461 29 463
rect 271 461 273 463
rect 291 460 293 462
rect 296 460 298 462
rect 33 458 35 460
rect 265 458 267 460
rect 2 455 4 457
rect 7 455 9 457
rect 27 456 29 458
rect 271 456 273 458
rect 291 455 293 457
rect 296 455 298 457
rect 2 450 4 452
rect 7 450 9 452
rect 27 451 29 453
rect 271 451 273 453
rect 291 450 293 452
rect 296 450 298 452
rect 2 445 4 447
rect 7 445 9 447
rect 27 446 29 448
rect 42 446 44 448
rect 47 446 49 448
rect 52 446 54 448
rect 57 446 59 448
rect 62 446 64 448
rect 67 446 69 448
rect 72 446 74 448
rect 77 446 79 448
rect 82 446 84 448
rect 87 446 89 448
rect 92 446 94 448
rect 97 446 99 448
rect 102 446 104 448
rect 107 446 109 448
rect 112 446 114 448
rect 117 446 119 448
rect 181 446 183 448
rect 186 446 188 448
rect 191 446 193 448
rect 196 446 198 448
rect 201 446 203 448
rect 206 446 208 448
rect 211 446 213 448
rect 216 446 218 448
rect 221 446 223 448
rect 226 446 228 448
rect 231 446 233 448
rect 236 446 238 448
rect 241 446 243 448
rect 246 446 248 448
rect 251 446 253 448
rect 256 446 258 448
rect 271 446 273 448
rect 291 445 293 447
rect 296 445 298 447
rect 2 440 4 442
rect 7 440 9 442
rect 291 440 293 442
rect 296 440 298 442
rect 22 438 24 440
rect 27 438 29 440
rect 32 438 34 440
rect 37 438 39 440
rect 42 438 44 440
rect 47 438 49 440
rect 52 438 54 440
rect 57 438 59 440
rect 62 438 64 440
rect 67 438 69 440
rect 72 438 74 440
rect 77 438 79 440
rect 82 438 84 440
rect 87 438 89 440
rect 92 438 94 440
rect 97 438 99 440
rect 102 438 104 440
rect 107 438 109 440
rect 112 438 114 440
rect 117 438 119 440
rect 181 438 183 440
rect 186 438 188 440
rect 191 438 193 440
rect 196 438 198 440
rect 201 438 203 440
rect 206 438 208 440
rect 211 438 213 440
rect 216 438 218 440
rect 221 438 223 440
rect 226 438 228 440
rect 231 438 233 440
rect 236 438 238 440
rect 241 438 243 440
rect 246 438 248 440
rect 251 438 253 440
rect 256 438 258 440
rect 261 438 263 440
rect 266 438 268 440
rect 271 438 273 440
rect 276 438 278 440
rect 2 435 4 437
rect 7 435 9 437
rect 291 435 293 437
rect 296 435 298 437
rect 22 433 24 435
rect 27 433 29 435
rect 32 433 34 435
rect 37 433 39 435
rect 42 433 44 435
rect 47 433 49 435
rect 52 433 54 435
rect 57 433 59 435
rect 62 433 64 435
rect 67 433 69 435
rect 72 433 74 435
rect 77 433 79 435
rect 82 433 84 435
rect 87 433 89 435
rect 92 433 94 435
rect 97 433 99 435
rect 102 433 104 435
rect 107 433 109 435
rect 112 433 114 435
rect 117 433 119 435
rect 181 433 183 435
rect 186 433 188 435
rect 191 433 193 435
rect 196 433 198 435
rect 201 433 203 435
rect 206 433 208 435
rect 211 433 213 435
rect 216 433 218 435
rect 221 433 223 435
rect 226 433 228 435
rect 231 433 233 435
rect 236 433 238 435
rect 241 433 243 435
rect 246 433 248 435
rect 251 433 253 435
rect 256 433 258 435
rect 261 433 263 435
rect 266 433 268 435
rect 271 433 273 435
rect 276 433 278 435
rect 2 430 4 432
rect 7 430 9 432
rect 291 430 293 432
rect 296 430 298 432
rect 2 425 4 427
rect 7 425 9 427
rect 291 425 293 427
rect 296 425 298 427
rect 4 415 6 417
rect 9 415 11 417
rect 14 415 16 417
rect 19 415 21 417
rect 24 415 26 417
rect 29 415 31 417
rect 34 415 36 417
rect 39 415 41 417
rect 44 415 46 417
rect 49 415 51 417
rect 54 415 56 417
rect 59 415 61 417
rect 64 415 66 417
rect 69 415 71 417
rect 74 415 76 417
rect 79 415 81 417
rect 84 415 86 417
rect 89 415 91 417
rect 94 415 96 417
rect 99 415 101 417
rect 104 415 106 417
rect 109 415 111 417
rect 114 415 116 417
rect 119 415 121 417
rect 124 415 126 417
rect 129 415 131 417
rect 134 415 136 417
rect 139 415 141 417
rect 144 415 146 417
rect 149 415 151 417
rect 154 415 156 417
rect 159 415 161 417
rect 164 415 166 417
rect 169 415 171 417
rect 174 415 176 417
rect 179 415 181 417
rect 184 415 186 417
rect 189 415 191 417
rect 194 415 196 417
rect 199 415 201 417
rect 204 415 206 417
rect 209 415 211 417
rect 214 415 216 417
rect 219 415 221 417
rect 224 415 226 417
rect 229 415 231 417
rect 234 415 236 417
rect 239 415 241 417
rect 244 415 246 417
rect 249 415 251 417
rect 254 415 256 417
rect 259 415 261 417
rect 264 415 266 417
rect 269 415 271 417
rect 274 415 276 417
rect 279 415 281 417
rect 284 415 286 417
rect 289 415 291 417
rect 294 415 296 417
rect 4 405 6 407
rect 9 405 11 407
rect 14 405 16 407
rect 19 405 21 407
rect 24 405 26 407
rect 29 405 31 407
rect 34 405 36 407
rect 39 405 41 407
rect 44 405 46 407
rect 49 405 51 407
rect 54 405 56 407
rect 59 405 61 407
rect 64 405 66 407
rect 69 405 71 407
rect 74 405 76 407
rect 79 405 81 407
rect 84 405 86 407
rect 89 405 91 407
rect 94 405 96 407
rect 99 405 101 407
rect 104 405 106 407
rect 109 405 111 407
rect 114 405 116 407
rect 119 405 121 407
rect 124 405 126 407
rect 129 405 131 407
rect 134 405 136 407
rect 139 405 141 407
rect 144 405 146 407
rect 149 405 151 407
rect 154 405 156 407
rect 159 405 161 407
rect 164 405 166 407
rect 169 405 171 407
rect 174 405 176 407
rect 179 405 181 407
rect 184 405 186 407
rect 189 405 191 407
rect 194 405 196 407
rect 199 405 201 407
rect 204 405 206 407
rect 209 405 211 407
rect 214 405 216 407
rect 219 405 221 407
rect 224 405 226 407
rect 229 405 231 407
rect 234 405 236 407
rect 239 405 241 407
rect 244 405 246 407
rect 249 405 251 407
rect 254 405 256 407
rect 259 405 261 407
rect 264 405 266 407
rect 269 405 271 407
rect 274 405 276 407
rect 279 405 281 407
rect 284 405 286 407
rect 289 405 291 407
rect 294 405 296 407
rect 4 395 6 397
rect 9 395 11 397
rect 14 395 16 397
rect 19 395 21 397
rect 24 395 26 397
rect 29 395 31 397
rect 34 395 36 397
rect 39 395 41 397
rect 44 395 46 397
rect 49 395 51 397
rect 54 395 56 397
rect 59 395 61 397
rect 64 395 66 397
rect 69 395 71 397
rect 74 395 76 397
rect 79 395 81 397
rect 84 395 86 397
rect 89 395 91 397
rect 94 395 96 397
rect 99 395 101 397
rect 104 395 106 397
rect 109 395 111 397
rect 114 395 116 397
rect 119 395 121 397
rect 124 395 126 397
rect 129 395 131 397
rect 134 395 136 397
rect 139 395 141 397
rect 144 395 146 397
rect 149 395 151 397
rect 154 395 156 397
rect 159 395 161 397
rect 164 395 166 397
rect 169 395 171 397
rect 174 395 176 397
rect 179 395 181 397
rect 184 395 186 397
rect 189 395 191 397
rect 194 395 196 397
rect 199 395 201 397
rect 204 395 206 397
rect 209 395 211 397
rect 214 395 216 397
rect 219 395 221 397
rect 224 395 226 397
rect 229 395 231 397
rect 234 395 236 397
rect 239 395 241 397
rect 244 395 246 397
rect 249 395 251 397
rect 254 395 256 397
rect 259 395 261 397
rect 264 395 266 397
rect 269 395 271 397
rect 274 395 276 397
rect 279 395 281 397
rect 284 395 286 397
rect 289 395 291 397
rect 294 395 296 397
rect 4 385 6 387
rect 9 385 11 387
rect 14 385 16 387
rect 19 385 21 387
rect 24 385 26 387
rect 29 385 31 387
rect 34 385 36 387
rect 39 385 41 387
rect 44 385 46 387
rect 49 385 51 387
rect 54 385 56 387
rect 59 385 61 387
rect 64 385 66 387
rect 69 385 71 387
rect 74 385 76 387
rect 79 385 81 387
rect 84 385 86 387
rect 89 385 91 387
rect 94 385 96 387
rect 99 385 101 387
rect 104 385 106 387
rect 109 385 111 387
rect 114 385 116 387
rect 119 385 121 387
rect 124 385 126 387
rect 129 385 131 387
rect 134 385 136 387
rect 139 385 141 387
rect 144 385 146 387
rect 149 385 151 387
rect 154 385 156 387
rect 159 385 161 387
rect 164 385 166 387
rect 169 385 171 387
rect 174 385 176 387
rect 179 385 181 387
rect 184 385 186 387
rect 189 385 191 387
rect 194 385 196 387
rect 199 385 201 387
rect 204 385 206 387
rect 209 385 211 387
rect 214 385 216 387
rect 219 385 221 387
rect 224 385 226 387
rect 229 385 231 387
rect 234 385 236 387
rect 239 385 241 387
rect 244 385 246 387
rect 249 385 251 387
rect 254 385 256 387
rect 259 385 261 387
rect 264 385 266 387
rect 269 385 271 387
rect 274 385 276 387
rect 279 385 281 387
rect 284 385 286 387
rect 289 385 291 387
rect 294 385 296 387
rect 4 375 6 377
rect 9 375 11 377
rect 14 375 16 377
rect 19 375 21 377
rect 24 375 26 377
rect 29 375 31 377
rect 34 375 36 377
rect 39 375 41 377
rect 44 375 46 377
rect 49 375 51 377
rect 54 375 56 377
rect 59 375 61 377
rect 64 375 66 377
rect 69 375 71 377
rect 74 375 76 377
rect 79 375 81 377
rect 84 375 86 377
rect 89 375 91 377
rect 94 375 96 377
rect 99 375 101 377
rect 104 375 106 377
rect 109 375 111 377
rect 114 375 116 377
rect 119 375 121 377
rect 124 375 126 377
rect 129 375 131 377
rect 134 375 136 377
rect 139 375 141 377
rect 144 375 146 377
rect 149 375 151 377
rect 154 375 156 377
rect 159 375 161 377
rect 164 375 166 377
rect 169 375 171 377
rect 174 375 176 377
rect 179 375 181 377
rect 184 375 186 377
rect 189 375 191 377
rect 194 375 196 377
rect 199 375 201 377
rect 204 375 206 377
rect 209 375 211 377
rect 214 375 216 377
rect 219 375 221 377
rect 224 375 226 377
rect 229 375 231 377
rect 234 375 236 377
rect 239 375 241 377
rect 244 375 246 377
rect 249 375 251 377
rect 254 375 256 377
rect 259 375 261 377
rect 264 375 266 377
rect 269 375 271 377
rect 274 375 276 377
rect 279 375 281 377
rect 284 375 286 377
rect 289 375 291 377
rect 294 375 296 377
rect 4 365 6 367
rect 9 365 11 367
rect 14 365 16 367
rect 19 365 21 367
rect 24 365 26 367
rect 29 365 31 367
rect 34 365 36 367
rect 39 365 41 367
rect 44 365 46 367
rect 49 365 51 367
rect 54 365 56 367
rect 59 365 61 367
rect 64 365 66 367
rect 69 365 71 367
rect 74 365 76 367
rect 79 365 81 367
rect 84 365 86 367
rect 89 365 91 367
rect 94 365 96 367
rect 99 365 101 367
rect 104 365 106 367
rect 109 365 111 367
rect 114 365 116 367
rect 119 365 121 367
rect 124 365 126 367
rect 129 365 131 367
rect 134 365 136 367
rect 139 365 141 367
rect 144 365 146 367
rect 149 365 151 367
rect 154 365 156 367
rect 159 365 161 367
rect 164 365 166 367
rect 169 365 171 367
rect 174 365 176 367
rect 179 365 181 367
rect 184 365 186 367
rect 189 365 191 367
rect 194 365 196 367
rect 199 365 201 367
rect 204 365 206 367
rect 209 365 211 367
rect 214 365 216 367
rect 219 365 221 367
rect 224 365 226 367
rect 229 365 231 367
rect 234 365 236 367
rect 239 365 241 367
rect 244 365 246 367
rect 249 365 251 367
rect 254 365 256 367
rect 259 365 261 367
rect 264 365 266 367
rect 269 365 271 367
rect 274 365 276 367
rect 279 365 281 367
rect 284 365 286 367
rect 289 365 291 367
rect 294 365 296 367
rect 4 355 6 357
rect 9 355 11 357
rect 14 355 16 357
rect 19 355 21 357
rect 24 355 26 357
rect 29 355 31 357
rect 34 355 36 357
rect 39 355 41 357
rect 44 355 46 357
rect 49 355 51 357
rect 54 355 56 357
rect 59 355 61 357
rect 64 355 66 357
rect 69 355 71 357
rect 74 355 76 357
rect 79 355 81 357
rect 84 355 86 357
rect 89 355 91 357
rect 94 355 96 357
rect 99 355 101 357
rect 104 355 106 357
rect 109 355 111 357
rect 114 355 116 357
rect 119 355 121 357
rect 124 355 126 357
rect 129 355 131 357
rect 134 355 136 357
rect 139 355 141 357
rect 144 355 146 357
rect 149 355 151 357
rect 154 355 156 357
rect 159 355 161 357
rect 164 355 166 357
rect 169 355 171 357
rect 174 355 176 357
rect 179 355 181 357
rect 184 355 186 357
rect 189 355 191 357
rect 194 355 196 357
rect 199 355 201 357
rect 204 355 206 357
rect 209 355 211 357
rect 214 355 216 357
rect 219 355 221 357
rect 224 355 226 357
rect 229 355 231 357
rect 234 355 236 357
rect 239 355 241 357
rect 244 355 246 357
rect 249 355 251 357
rect 254 355 256 357
rect 259 355 261 357
rect 264 355 266 357
rect 269 355 271 357
rect 274 355 276 357
rect 279 355 281 357
rect 284 355 286 357
rect 289 355 291 357
rect 294 355 296 357
rect 4 345 6 347
rect 9 345 11 347
rect 14 345 16 347
rect 19 345 21 347
rect 24 345 26 347
rect 29 345 31 347
rect 34 345 36 347
rect 39 345 41 347
rect 44 345 46 347
rect 49 345 51 347
rect 54 345 56 347
rect 59 345 61 347
rect 64 345 66 347
rect 69 345 71 347
rect 74 345 76 347
rect 79 345 81 347
rect 84 345 86 347
rect 89 345 91 347
rect 94 345 96 347
rect 99 345 101 347
rect 104 345 106 347
rect 109 345 111 347
rect 114 345 116 347
rect 119 345 121 347
rect 124 345 126 347
rect 129 345 131 347
rect 134 345 136 347
rect 139 345 141 347
rect 144 345 146 347
rect 149 345 151 347
rect 154 345 156 347
rect 159 345 161 347
rect 164 345 166 347
rect 169 345 171 347
rect 174 345 176 347
rect 179 345 181 347
rect 184 345 186 347
rect 189 345 191 347
rect 194 345 196 347
rect 199 345 201 347
rect 204 345 206 347
rect 209 345 211 347
rect 214 345 216 347
rect 219 345 221 347
rect 224 345 226 347
rect 229 345 231 347
rect 234 345 236 347
rect 239 345 241 347
rect 244 345 246 347
rect 249 345 251 347
rect 254 345 256 347
rect 259 345 261 347
rect 264 345 266 347
rect 269 345 271 347
rect 274 345 276 347
rect 279 345 281 347
rect 284 345 286 347
rect 289 345 291 347
rect 294 345 296 347
rect 3 323 5 325
rect 8 323 10 325
rect 13 323 15 325
rect 18 323 20 325
rect 23 323 25 325
rect 28 323 30 325
rect 33 323 35 325
rect 38 323 40 325
rect 43 323 45 325
rect 48 323 50 325
rect 53 323 55 325
rect 58 323 60 325
rect 63 323 65 325
rect 68 323 70 325
rect 73 323 75 325
rect 78 323 80 325
rect 83 323 85 325
rect 88 323 90 325
rect 93 323 95 325
rect 144 323 146 325
rect 149 323 151 325
rect 154 323 156 325
rect 205 323 207 325
rect 210 323 212 325
rect 215 323 217 325
rect 220 323 222 325
rect 225 323 227 325
rect 230 323 232 325
rect 235 323 237 325
rect 240 323 242 325
rect 245 323 247 325
rect 250 323 252 325
rect 255 323 257 325
rect 260 323 262 325
rect 265 323 267 325
rect 270 323 272 325
rect 275 323 277 325
rect 280 323 282 325
rect 285 323 287 325
rect 290 323 292 325
rect 295 323 297 325
rect 3 313 5 315
rect 8 313 10 315
rect 13 313 15 315
rect 18 313 20 315
rect 23 313 25 315
rect 28 313 30 315
rect 33 313 35 315
rect 38 313 40 315
rect 43 313 45 315
rect 48 313 50 315
rect 53 313 55 315
rect 58 313 60 315
rect 63 313 65 315
rect 68 313 70 315
rect 73 313 75 315
rect 78 313 80 315
rect 83 313 85 315
rect 88 313 90 315
rect 93 313 95 315
rect 144 313 146 315
rect 149 313 151 315
rect 154 313 156 315
rect 205 313 207 315
rect 210 313 212 315
rect 215 313 217 315
rect 220 313 222 315
rect 225 313 227 315
rect 230 313 232 315
rect 235 313 237 315
rect 240 313 242 315
rect 245 313 247 315
rect 250 313 252 315
rect 255 313 257 315
rect 260 313 262 315
rect 265 313 267 315
rect 270 313 272 315
rect 275 313 277 315
rect 280 313 282 315
rect 285 313 287 315
rect 290 313 292 315
rect 295 313 297 315
rect 3 303 5 305
rect 8 303 10 305
rect 13 303 15 305
rect 18 303 20 305
rect 23 303 25 305
rect 28 303 30 305
rect 33 303 35 305
rect 38 303 40 305
rect 43 303 45 305
rect 48 303 50 305
rect 53 303 55 305
rect 58 303 60 305
rect 63 303 65 305
rect 68 303 70 305
rect 73 303 75 305
rect 78 303 80 305
rect 83 303 85 305
rect 88 303 90 305
rect 93 303 95 305
rect 144 303 146 305
rect 149 303 151 305
rect 154 303 156 305
rect 205 303 207 305
rect 210 303 212 305
rect 215 303 217 305
rect 220 303 222 305
rect 225 303 227 305
rect 230 303 232 305
rect 235 303 237 305
rect 240 303 242 305
rect 245 303 247 305
rect 250 303 252 305
rect 255 303 257 305
rect 260 303 262 305
rect 265 303 267 305
rect 270 303 272 305
rect 275 303 277 305
rect 280 303 282 305
rect 285 303 287 305
rect 290 303 292 305
rect 295 303 297 305
rect 3 293 5 295
rect 8 293 10 295
rect 13 293 15 295
rect 18 293 20 295
rect 23 293 25 295
rect 28 293 30 295
rect 33 293 35 295
rect 38 293 40 295
rect 43 293 45 295
rect 48 293 50 295
rect 53 293 55 295
rect 58 293 60 295
rect 63 293 65 295
rect 68 293 70 295
rect 73 293 75 295
rect 78 293 80 295
rect 83 293 85 295
rect 88 293 90 295
rect 93 293 95 295
rect 144 293 146 295
rect 149 293 151 295
rect 154 293 156 295
rect 205 293 207 295
rect 210 293 212 295
rect 215 293 217 295
rect 220 293 222 295
rect 225 293 227 295
rect 230 293 232 295
rect 235 293 237 295
rect 240 293 242 295
rect 245 293 247 295
rect 250 293 252 295
rect 255 293 257 295
rect 260 293 262 295
rect 265 293 267 295
rect 270 293 272 295
rect 275 293 277 295
rect 280 293 282 295
rect 285 293 287 295
rect 290 293 292 295
rect 295 293 297 295
rect 3 283 5 285
rect 8 283 10 285
rect 13 283 15 285
rect 18 283 20 285
rect 23 283 25 285
rect 28 283 30 285
rect 33 283 35 285
rect 38 283 40 285
rect 43 283 45 285
rect 48 283 50 285
rect 53 283 55 285
rect 58 283 60 285
rect 63 283 65 285
rect 68 283 70 285
rect 73 283 75 285
rect 78 283 80 285
rect 83 283 85 285
rect 88 283 90 285
rect 93 283 95 285
rect 144 283 146 285
rect 149 283 151 285
rect 154 283 156 285
rect 205 283 207 285
rect 210 283 212 285
rect 215 283 217 285
rect 220 283 222 285
rect 225 283 227 285
rect 230 283 232 285
rect 235 283 237 285
rect 240 283 242 285
rect 245 283 247 285
rect 250 283 252 285
rect 255 283 257 285
rect 260 283 262 285
rect 265 283 267 285
rect 270 283 272 285
rect 275 283 277 285
rect 280 283 282 285
rect 285 283 287 285
rect 290 283 292 285
rect 295 283 297 285
rect 3 273 5 275
rect 8 273 10 275
rect 13 273 15 275
rect 18 273 20 275
rect 23 273 25 275
rect 28 273 30 275
rect 33 273 35 275
rect 38 273 40 275
rect 43 273 45 275
rect 48 273 50 275
rect 53 273 55 275
rect 58 273 60 275
rect 63 273 65 275
rect 68 273 70 275
rect 73 273 75 275
rect 78 273 80 275
rect 83 273 85 275
rect 88 273 90 275
rect 93 273 95 275
rect 144 273 146 275
rect 149 273 151 275
rect 154 273 156 275
rect 205 273 207 275
rect 210 273 212 275
rect 215 273 217 275
rect 220 273 222 275
rect 225 273 227 275
rect 230 273 232 275
rect 235 273 237 275
rect 240 273 242 275
rect 245 273 247 275
rect 250 273 252 275
rect 255 273 257 275
rect 260 273 262 275
rect 265 273 267 275
rect 270 273 272 275
rect 275 273 277 275
rect 280 273 282 275
rect 285 273 287 275
rect 290 273 292 275
rect 295 273 297 275
rect 3 263 5 265
rect 8 263 10 265
rect 13 263 15 265
rect 18 263 20 265
rect 23 263 25 265
rect 28 263 30 265
rect 33 263 35 265
rect 38 263 40 265
rect 43 263 45 265
rect 48 263 50 265
rect 53 263 55 265
rect 58 263 60 265
rect 63 263 65 265
rect 68 263 70 265
rect 73 263 75 265
rect 78 263 80 265
rect 83 263 85 265
rect 88 263 90 265
rect 93 263 95 265
rect 144 263 146 265
rect 149 263 151 265
rect 154 263 156 265
rect 205 263 207 265
rect 210 263 212 265
rect 215 263 217 265
rect 220 263 222 265
rect 225 263 227 265
rect 230 263 232 265
rect 235 263 237 265
rect 240 263 242 265
rect 245 263 247 265
rect 250 263 252 265
rect 255 263 257 265
rect 260 263 262 265
rect 265 263 267 265
rect 270 263 272 265
rect 275 263 277 265
rect 280 263 282 265
rect 285 263 287 265
rect 290 263 292 265
rect 295 263 297 265
rect 3 253 5 255
rect 9 253 11 255
rect 14 253 16 255
rect 19 253 21 255
rect 24 253 26 255
rect 29 253 31 255
rect 34 253 36 255
rect 39 253 41 255
rect 44 253 46 255
rect 49 253 51 255
rect 54 253 56 255
rect 59 253 61 255
rect 64 253 66 255
rect 69 253 71 255
rect 74 253 76 255
rect 79 253 81 255
rect 84 253 86 255
rect 89 253 91 255
rect 94 253 96 255
rect 144 253 146 255
rect 149 253 151 255
rect 154 253 156 255
rect 204 253 206 255
rect 209 253 211 255
rect 214 253 216 255
rect 219 253 221 255
rect 224 253 226 255
rect 229 253 231 255
rect 234 253 236 255
rect 239 253 241 255
rect 244 253 246 255
rect 249 253 251 255
rect 254 253 256 255
rect 259 253 261 255
rect 264 253 266 255
rect 269 253 271 255
rect 274 253 276 255
rect 279 253 281 255
rect 284 253 286 255
rect 289 253 291 255
rect 295 253 297 255
rect 3 248 5 250
rect 295 248 297 250
rect 3 243 5 245
rect 16 242 18 244
rect 21 242 23 244
rect 26 242 28 244
rect 31 242 33 244
rect 36 242 38 244
rect 41 242 43 244
rect 46 242 48 244
rect 51 242 53 244
rect 56 242 58 244
rect 61 242 63 244
rect 66 242 68 244
rect 71 242 73 244
rect 76 242 78 244
rect 81 242 83 244
rect 86 242 88 244
rect 91 242 93 244
rect 96 242 98 244
rect 101 242 103 244
rect 106 242 108 244
rect 111 242 113 244
rect 116 242 118 244
rect 121 242 123 244
rect 126 242 128 244
rect 131 242 133 244
rect 136 242 138 244
rect 141 242 143 244
rect 146 242 148 244
rect 151 242 153 244
rect 156 242 158 244
rect 161 242 163 244
rect 166 242 168 244
rect 171 242 173 244
rect 176 242 178 244
rect 181 242 183 244
rect 186 242 188 244
rect 191 242 193 244
rect 196 242 198 244
rect 201 242 203 244
rect 206 242 208 244
rect 211 242 213 244
rect 216 242 218 244
rect 221 242 223 244
rect 226 242 228 244
rect 231 242 233 244
rect 236 242 238 244
rect 241 242 243 244
rect 246 242 248 244
rect 251 242 253 244
rect 256 242 258 244
rect 261 242 263 244
rect 266 242 268 244
rect 271 242 273 244
rect 276 242 278 244
rect 281 242 283 244
rect 295 243 297 245
rect 3 238 5 240
rect 16 237 18 239
rect 21 237 23 239
rect 26 237 28 239
rect 31 237 33 239
rect 36 237 38 239
rect 41 237 43 239
rect 46 237 48 239
rect 51 237 53 239
rect 56 237 58 239
rect 61 237 63 239
rect 66 237 68 239
rect 71 237 73 239
rect 76 237 78 239
rect 81 237 83 239
rect 86 237 88 239
rect 91 237 93 239
rect 96 237 98 239
rect 101 237 103 239
rect 106 237 108 239
rect 111 237 113 239
rect 116 237 118 239
rect 121 237 123 239
rect 126 237 128 239
rect 131 237 133 239
rect 136 237 138 239
rect 141 237 143 239
rect 146 237 148 239
rect 151 237 153 239
rect 156 237 158 239
rect 161 237 163 239
rect 166 237 168 239
rect 171 237 173 239
rect 176 237 178 239
rect 181 237 183 239
rect 186 237 188 239
rect 191 237 193 239
rect 196 237 198 239
rect 201 237 203 239
rect 206 237 208 239
rect 211 237 213 239
rect 216 237 218 239
rect 221 237 223 239
rect 226 237 228 239
rect 231 237 233 239
rect 236 237 238 239
rect 241 237 243 239
rect 246 237 248 239
rect 251 237 253 239
rect 256 237 258 239
rect 261 237 263 239
rect 266 237 268 239
rect 271 237 273 239
rect 276 237 278 239
rect 281 237 283 239
rect 295 238 297 240
rect 3 233 5 235
rect 16 232 18 234
rect 21 232 23 234
rect 26 232 28 234
rect 31 232 33 234
rect 36 232 38 234
rect 41 232 43 234
rect 46 232 48 234
rect 51 232 53 234
rect 56 232 58 234
rect 61 232 63 234
rect 66 232 68 234
rect 71 232 73 234
rect 76 232 78 234
rect 81 232 83 234
rect 86 232 88 234
rect 91 232 93 234
rect 96 232 98 234
rect 101 232 103 234
rect 106 232 108 234
rect 111 232 113 234
rect 116 232 118 234
rect 121 232 123 234
rect 126 232 128 234
rect 131 232 133 234
rect 136 232 138 234
rect 141 232 143 234
rect 146 232 148 234
rect 151 232 153 234
rect 156 232 158 234
rect 161 232 163 234
rect 166 232 168 234
rect 171 232 173 234
rect 176 232 178 234
rect 181 232 183 234
rect 186 232 188 234
rect 191 232 193 234
rect 196 232 198 234
rect 201 232 203 234
rect 206 232 208 234
rect 211 232 213 234
rect 216 232 218 234
rect 221 232 223 234
rect 226 232 228 234
rect 231 232 233 234
rect 236 232 238 234
rect 241 232 243 234
rect 246 232 248 234
rect 251 232 253 234
rect 256 232 258 234
rect 261 232 263 234
rect 266 232 268 234
rect 271 232 273 234
rect 276 232 278 234
rect 281 232 283 234
rect 295 233 297 235
rect 3 228 5 230
rect 295 228 297 230
rect 16 226 18 228
rect 21 226 23 228
rect 26 226 28 228
rect 31 226 33 228
rect 36 226 38 228
rect 41 226 43 228
rect 46 226 48 228
rect 51 226 53 228
rect 56 226 58 228
rect 61 226 63 228
rect 66 226 68 228
rect 71 226 73 228
rect 76 226 78 228
rect 81 226 83 228
rect 86 226 88 228
rect 91 226 93 228
rect 96 226 98 228
rect 101 226 103 228
rect 106 226 108 228
rect 111 226 113 228
rect 116 226 118 228
rect 121 226 123 228
rect 126 226 128 228
rect 131 226 133 228
rect 136 226 138 228
rect 141 226 143 228
rect 146 226 148 228
rect 151 226 153 228
rect 156 226 158 228
rect 161 226 163 228
rect 166 226 168 228
rect 171 226 173 228
rect 176 226 178 228
rect 181 226 183 228
rect 186 226 188 228
rect 191 226 193 228
rect 196 226 198 228
rect 201 226 203 228
rect 206 226 208 228
rect 211 226 213 228
rect 216 226 218 228
rect 221 226 223 228
rect 226 226 228 228
rect 231 226 233 228
rect 236 226 238 228
rect 241 226 243 228
rect 246 226 248 228
rect 251 226 253 228
rect 256 226 258 228
rect 261 226 263 228
rect 266 226 268 228
rect 271 226 273 228
rect 276 226 278 228
rect 281 226 283 228
rect 3 223 5 225
rect 295 223 297 225
rect 3 218 5 220
rect 295 218 297 220
rect 16 216 18 218
rect 21 216 23 218
rect 26 216 28 218
rect 31 216 33 218
rect 36 216 38 218
rect 41 216 43 218
rect 46 216 48 218
rect 51 216 53 218
rect 56 216 58 218
rect 61 216 63 218
rect 66 216 68 218
rect 71 216 73 218
rect 76 216 78 218
rect 81 216 83 218
rect 86 216 88 218
rect 91 216 93 218
rect 96 216 98 218
rect 101 216 103 218
rect 106 216 108 218
rect 111 216 113 218
rect 116 216 118 218
rect 121 216 123 218
rect 126 216 128 218
rect 131 216 133 218
rect 136 216 138 218
rect 141 216 143 218
rect 146 216 148 218
rect 151 216 153 218
rect 156 216 158 218
rect 161 216 163 218
rect 166 216 168 218
rect 171 216 173 218
rect 176 216 178 218
rect 181 216 183 218
rect 186 216 188 218
rect 191 216 193 218
rect 196 216 198 218
rect 201 216 203 218
rect 206 216 208 218
rect 211 216 213 218
rect 216 216 218 218
rect 221 216 223 218
rect 226 216 228 218
rect 231 216 233 218
rect 236 216 238 218
rect 241 216 243 218
rect 246 216 248 218
rect 251 216 253 218
rect 256 216 258 218
rect 261 216 263 218
rect 266 216 268 218
rect 271 216 273 218
rect 276 216 278 218
rect 281 216 283 218
rect 3 213 5 215
rect 295 213 297 215
rect 3 208 5 210
rect 295 208 297 210
rect 16 206 18 208
rect 21 206 23 208
rect 26 206 28 208
rect 31 206 33 208
rect 36 206 38 208
rect 41 206 43 208
rect 46 206 48 208
rect 51 206 53 208
rect 56 206 58 208
rect 61 206 63 208
rect 66 206 68 208
rect 71 206 73 208
rect 76 206 78 208
rect 81 206 83 208
rect 86 206 88 208
rect 91 206 93 208
rect 96 206 98 208
rect 101 206 103 208
rect 106 206 108 208
rect 111 206 113 208
rect 116 206 118 208
rect 121 206 123 208
rect 126 206 128 208
rect 131 206 133 208
rect 136 206 138 208
rect 141 206 143 208
rect 146 206 148 208
rect 151 206 153 208
rect 156 206 158 208
rect 161 206 163 208
rect 166 206 168 208
rect 171 206 173 208
rect 176 206 178 208
rect 181 206 183 208
rect 186 206 188 208
rect 191 206 193 208
rect 196 206 198 208
rect 201 206 203 208
rect 206 206 208 208
rect 211 206 213 208
rect 216 206 218 208
rect 221 206 223 208
rect 226 206 228 208
rect 231 206 233 208
rect 236 206 238 208
rect 241 206 243 208
rect 246 206 248 208
rect 251 206 253 208
rect 256 206 258 208
rect 261 206 263 208
rect 266 206 268 208
rect 271 206 273 208
rect 276 206 278 208
rect 281 206 283 208
rect 3 203 5 205
rect 295 203 297 205
rect 3 198 5 200
rect 295 198 297 200
rect 16 196 18 198
rect 21 196 23 198
rect 26 196 28 198
rect 31 196 33 198
rect 36 196 38 198
rect 41 196 43 198
rect 46 196 48 198
rect 51 196 53 198
rect 56 196 58 198
rect 61 196 63 198
rect 66 196 68 198
rect 71 196 73 198
rect 76 196 78 198
rect 81 196 83 198
rect 86 196 88 198
rect 91 196 93 198
rect 96 196 98 198
rect 101 196 103 198
rect 106 196 108 198
rect 111 196 113 198
rect 116 196 118 198
rect 121 196 123 198
rect 126 196 128 198
rect 131 196 133 198
rect 136 196 138 198
rect 141 196 143 198
rect 146 196 148 198
rect 151 196 153 198
rect 156 196 158 198
rect 161 196 163 198
rect 166 196 168 198
rect 171 196 173 198
rect 176 196 178 198
rect 181 196 183 198
rect 186 196 188 198
rect 191 196 193 198
rect 196 196 198 198
rect 201 196 203 198
rect 206 196 208 198
rect 211 196 213 198
rect 216 196 218 198
rect 221 196 223 198
rect 226 196 228 198
rect 231 196 233 198
rect 236 196 238 198
rect 241 196 243 198
rect 246 196 248 198
rect 251 196 253 198
rect 256 196 258 198
rect 261 196 263 198
rect 266 196 268 198
rect 271 196 273 198
rect 276 196 278 198
rect 281 196 283 198
rect 3 193 5 195
rect 295 193 297 195
rect 3 188 5 190
rect 295 188 297 190
rect 16 186 18 188
rect 21 186 23 188
rect 26 186 28 188
rect 31 186 33 188
rect 36 186 38 188
rect 41 186 43 188
rect 46 186 48 188
rect 51 186 53 188
rect 56 186 58 188
rect 61 186 63 188
rect 66 186 68 188
rect 71 186 73 188
rect 76 186 78 188
rect 81 186 83 188
rect 86 186 88 188
rect 91 186 93 188
rect 96 186 98 188
rect 101 186 103 188
rect 106 186 108 188
rect 111 186 113 188
rect 116 186 118 188
rect 121 186 123 188
rect 126 186 128 188
rect 131 186 133 188
rect 136 186 138 188
rect 141 186 143 188
rect 146 186 148 188
rect 151 186 153 188
rect 156 186 158 188
rect 161 186 163 188
rect 166 186 168 188
rect 171 186 173 188
rect 176 186 178 188
rect 181 186 183 188
rect 186 186 188 188
rect 191 186 193 188
rect 196 186 198 188
rect 201 186 203 188
rect 206 186 208 188
rect 211 186 213 188
rect 216 186 218 188
rect 221 186 223 188
rect 226 186 228 188
rect 231 186 233 188
rect 236 186 238 188
rect 241 186 243 188
rect 246 186 248 188
rect 251 186 253 188
rect 256 186 258 188
rect 261 186 263 188
rect 266 186 268 188
rect 271 186 273 188
rect 276 186 278 188
rect 281 186 283 188
rect 3 183 5 185
rect 295 183 297 185
rect 3 178 5 180
rect 295 178 297 180
rect 16 176 18 178
rect 21 176 23 178
rect 26 176 28 178
rect 31 176 33 178
rect 36 176 38 178
rect 41 176 43 178
rect 46 176 48 178
rect 51 176 53 178
rect 56 176 58 178
rect 61 176 63 178
rect 66 176 68 178
rect 71 176 73 178
rect 76 176 78 178
rect 81 176 83 178
rect 86 176 88 178
rect 91 176 93 178
rect 96 176 98 178
rect 101 176 103 178
rect 106 176 108 178
rect 111 176 113 178
rect 116 176 118 178
rect 121 176 123 178
rect 126 176 128 178
rect 131 176 133 178
rect 136 176 138 178
rect 141 176 143 178
rect 146 176 148 178
rect 151 176 153 178
rect 156 176 158 178
rect 161 176 163 178
rect 166 176 168 178
rect 171 176 173 178
rect 176 176 178 178
rect 181 176 183 178
rect 186 176 188 178
rect 191 176 193 178
rect 196 176 198 178
rect 201 176 203 178
rect 206 176 208 178
rect 211 176 213 178
rect 216 176 218 178
rect 221 176 223 178
rect 226 176 228 178
rect 231 176 233 178
rect 236 176 238 178
rect 241 176 243 178
rect 246 176 248 178
rect 251 176 253 178
rect 256 176 258 178
rect 261 176 263 178
rect 266 176 268 178
rect 271 176 273 178
rect 276 176 278 178
rect 281 176 283 178
rect 3 173 5 175
rect 295 173 297 175
rect 3 168 5 170
rect 295 168 297 170
rect 16 166 18 168
rect 21 166 23 168
rect 26 166 28 168
rect 31 166 33 168
rect 36 166 38 168
rect 41 166 43 168
rect 46 166 48 168
rect 51 166 53 168
rect 56 166 58 168
rect 61 166 63 168
rect 66 166 68 168
rect 71 166 73 168
rect 76 166 78 168
rect 81 166 83 168
rect 86 166 88 168
rect 91 166 93 168
rect 96 166 98 168
rect 101 166 103 168
rect 106 166 108 168
rect 111 166 113 168
rect 116 166 118 168
rect 121 166 123 168
rect 126 166 128 168
rect 131 166 133 168
rect 136 166 138 168
rect 141 166 143 168
rect 146 166 148 168
rect 151 166 153 168
rect 156 166 158 168
rect 161 166 163 168
rect 166 166 168 168
rect 171 166 173 168
rect 176 166 178 168
rect 181 166 183 168
rect 186 166 188 168
rect 191 166 193 168
rect 196 166 198 168
rect 201 166 203 168
rect 206 166 208 168
rect 211 166 213 168
rect 216 166 218 168
rect 221 166 223 168
rect 226 166 228 168
rect 231 166 233 168
rect 236 166 238 168
rect 241 166 243 168
rect 246 166 248 168
rect 251 166 253 168
rect 256 166 258 168
rect 261 166 263 168
rect 266 166 268 168
rect 271 166 273 168
rect 276 166 278 168
rect 281 166 283 168
rect 3 163 5 165
rect 295 163 297 165
rect 3 158 5 160
rect 295 158 297 160
rect 16 156 18 158
rect 21 156 23 158
rect 26 156 28 158
rect 31 156 33 158
rect 36 156 38 158
rect 41 156 43 158
rect 46 156 48 158
rect 51 156 53 158
rect 56 156 58 158
rect 61 156 63 158
rect 66 156 68 158
rect 71 156 73 158
rect 76 156 78 158
rect 81 156 83 158
rect 86 156 88 158
rect 91 156 93 158
rect 96 156 98 158
rect 101 156 103 158
rect 106 156 108 158
rect 111 156 113 158
rect 116 156 118 158
rect 121 156 123 158
rect 126 156 128 158
rect 131 156 133 158
rect 136 156 138 158
rect 141 156 143 158
rect 146 156 148 158
rect 151 156 153 158
rect 156 156 158 158
rect 161 156 163 158
rect 166 156 168 158
rect 171 156 173 158
rect 176 156 178 158
rect 181 156 183 158
rect 186 156 188 158
rect 191 156 193 158
rect 196 156 198 158
rect 201 156 203 158
rect 206 156 208 158
rect 211 156 213 158
rect 216 156 218 158
rect 221 156 223 158
rect 226 156 228 158
rect 231 156 233 158
rect 236 156 238 158
rect 241 156 243 158
rect 246 156 248 158
rect 251 156 253 158
rect 256 156 258 158
rect 261 156 263 158
rect 266 156 268 158
rect 271 156 273 158
rect 276 156 278 158
rect 281 156 283 158
rect 3 153 5 155
rect 295 153 297 155
rect 3 148 5 150
rect 295 148 297 150
rect 16 146 18 148
rect 21 146 23 148
rect 26 146 28 148
rect 31 146 33 148
rect 36 146 38 148
rect 41 146 43 148
rect 46 146 48 148
rect 51 146 53 148
rect 56 146 58 148
rect 61 146 63 148
rect 66 146 68 148
rect 71 146 73 148
rect 76 146 78 148
rect 81 146 83 148
rect 86 146 88 148
rect 91 146 93 148
rect 96 146 98 148
rect 101 146 103 148
rect 106 146 108 148
rect 111 146 113 148
rect 116 146 118 148
rect 121 146 123 148
rect 126 146 128 148
rect 131 146 133 148
rect 136 146 138 148
rect 141 146 143 148
rect 146 146 148 148
rect 151 146 153 148
rect 156 146 158 148
rect 161 146 163 148
rect 166 146 168 148
rect 171 146 173 148
rect 176 146 178 148
rect 181 146 183 148
rect 186 146 188 148
rect 191 146 193 148
rect 196 146 198 148
rect 201 146 203 148
rect 206 146 208 148
rect 211 146 213 148
rect 216 146 218 148
rect 221 146 223 148
rect 226 146 228 148
rect 231 146 233 148
rect 236 146 238 148
rect 241 146 243 148
rect 246 146 248 148
rect 251 146 253 148
rect 256 146 258 148
rect 261 146 263 148
rect 266 146 268 148
rect 271 146 273 148
rect 276 146 278 148
rect 281 146 283 148
rect 3 143 5 145
rect 295 143 297 145
rect 3 138 5 140
rect 295 138 297 140
rect 16 136 18 138
rect 21 136 23 138
rect 26 136 28 138
rect 31 136 33 138
rect 36 136 38 138
rect 41 136 43 138
rect 46 136 48 138
rect 51 136 53 138
rect 56 136 58 138
rect 61 136 63 138
rect 66 136 68 138
rect 71 136 73 138
rect 76 136 78 138
rect 81 136 83 138
rect 86 136 88 138
rect 91 136 93 138
rect 96 136 98 138
rect 101 136 103 138
rect 106 136 108 138
rect 111 136 113 138
rect 116 136 118 138
rect 121 136 123 138
rect 126 136 128 138
rect 131 136 133 138
rect 136 136 138 138
rect 141 136 143 138
rect 146 136 148 138
rect 151 136 153 138
rect 156 136 158 138
rect 161 136 163 138
rect 166 136 168 138
rect 171 136 173 138
rect 176 136 178 138
rect 181 136 183 138
rect 186 136 188 138
rect 191 136 193 138
rect 196 136 198 138
rect 201 136 203 138
rect 206 136 208 138
rect 211 136 213 138
rect 216 136 218 138
rect 221 136 223 138
rect 226 136 228 138
rect 231 136 233 138
rect 236 136 238 138
rect 241 136 243 138
rect 246 136 248 138
rect 251 136 253 138
rect 256 136 258 138
rect 261 136 263 138
rect 266 136 268 138
rect 271 136 273 138
rect 276 136 278 138
rect 281 136 283 138
rect 3 133 5 135
rect 295 133 297 135
rect 3 128 5 130
rect 295 128 297 130
rect 16 126 18 128
rect 21 126 23 128
rect 26 126 28 128
rect 31 126 33 128
rect 36 126 38 128
rect 41 126 43 128
rect 46 126 48 128
rect 51 126 53 128
rect 56 126 58 128
rect 61 126 63 128
rect 66 126 68 128
rect 71 126 73 128
rect 76 126 78 128
rect 81 126 83 128
rect 86 126 88 128
rect 91 126 93 128
rect 96 126 98 128
rect 101 126 103 128
rect 106 126 108 128
rect 111 126 113 128
rect 116 126 118 128
rect 121 126 123 128
rect 126 126 128 128
rect 131 126 133 128
rect 136 126 138 128
rect 141 126 143 128
rect 146 126 148 128
rect 151 126 153 128
rect 156 126 158 128
rect 161 126 163 128
rect 166 126 168 128
rect 171 126 173 128
rect 176 126 178 128
rect 181 126 183 128
rect 186 126 188 128
rect 191 126 193 128
rect 196 126 198 128
rect 201 126 203 128
rect 206 126 208 128
rect 211 126 213 128
rect 216 126 218 128
rect 221 126 223 128
rect 226 126 228 128
rect 231 126 233 128
rect 236 126 238 128
rect 241 126 243 128
rect 246 126 248 128
rect 251 126 253 128
rect 256 126 258 128
rect 261 126 263 128
rect 266 126 268 128
rect 271 126 273 128
rect 276 126 278 128
rect 281 126 283 128
rect 3 123 5 125
rect 295 123 297 125
rect 3 118 5 120
rect 295 118 297 120
rect 16 116 18 118
rect 21 116 23 118
rect 26 116 28 118
rect 31 116 33 118
rect 36 116 38 118
rect 41 116 43 118
rect 46 116 48 118
rect 51 116 53 118
rect 56 116 58 118
rect 61 116 63 118
rect 66 116 68 118
rect 71 116 73 118
rect 76 116 78 118
rect 81 116 83 118
rect 86 116 88 118
rect 91 116 93 118
rect 96 116 98 118
rect 101 116 103 118
rect 106 116 108 118
rect 111 116 113 118
rect 116 116 118 118
rect 121 116 123 118
rect 126 116 128 118
rect 131 116 133 118
rect 136 116 138 118
rect 141 116 143 118
rect 146 116 148 118
rect 151 116 153 118
rect 156 116 158 118
rect 161 116 163 118
rect 166 116 168 118
rect 171 116 173 118
rect 176 116 178 118
rect 181 116 183 118
rect 186 116 188 118
rect 191 116 193 118
rect 196 116 198 118
rect 201 116 203 118
rect 206 116 208 118
rect 211 116 213 118
rect 216 116 218 118
rect 221 116 223 118
rect 226 116 228 118
rect 231 116 233 118
rect 236 116 238 118
rect 241 116 243 118
rect 246 116 248 118
rect 251 116 253 118
rect 256 116 258 118
rect 261 116 263 118
rect 266 116 268 118
rect 271 116 273 118
rect 276 116 278 118
rect 281 116 283 118
rect 3 113 5 115
rect 295 113 297 115
rect 3 108 5 110
rect 295 108 297 110
rect 16 106 18 108
rect 21 106 23 108
rect 26 106 28 108
rect 31 106 33 108
rect 36 106 38 108
rect 41 106 43 108
rect 46 106 48 108
rect 51 106 53 108
rect 56 106 58 108
rect 61 106 63 108
rect 66 106 68 108
rect 71 106 73 108
rect 76 106 78 108
rect 81 106 83 108
rect 86 106 88 108
rect 91 106 93 108
rect 96 106 98 108
rect 101 106 103 108
rect 106 106 108 108
rect 111 106 113 108
rect 116 106 118 108
rect 121 106 123 108
rect 126 106 128 108
rect 131 106 133 108
rect 136 106 138 108
rect 141 106 143 108
rect 146 106 148 108
rect 151 106 153 108
rect 156 106 158 108
rect 161 106 163 108
rect 166 106 168 108
rect 171 106 173 108
rect 176 106 178 108
rect 181 106 183 108
rect 186 106 188 108
rect 191 106 193 108
rect 196 106 198 108
rect 201 106 203 108
rect 206 106 208 108
rect 211 106 213 108
rect 216 106 218 108
rect 221 106 223 108
rect 226 106 228 108
rect 231 106 233 108
rect 236 106 238 108
rect 241 106 243 108
rect 246 106 248 108
rect 251 106 253 108
rect 256 106 258 108
rect 261 106 263 108
rect 266 106 268 108
rect 271 106 273 108
rect 276 106 278 108
rect 281 106 283 108
rect 3 103 5 105
rect 295 103 297 105
rect 3 98 5 100
rect 295 98 297 100
rect 16 96 18 98
rect 21 96 23 98
rect 26 96 28 98
rect 31 96 33 98
rect 36 96 38 98
rect 41 96 43 98
rect 46 96 48 98
rect 51 96 53 98
rect 56 96 58 98
rect 61 96 63 98
rect 66 96 68 98
rect 71 96 73 98
rect 76 96 78 98
rect 81 96 83 98
rect 86 96 88 98
rect 91 96 93 98
rect 96 96 98 98
rect 101 96 103 98
rect 106 96 108 98
rect 111 96 113 98
rect 116 96 118 98
rect 121 96 123 98
rect 126 96 128 98
rect 131 96 133 98
rect 136 96 138 98
rect 141 96 143 98
rect 146 96 148 98
rect 151 96 153 98
rect 156 96 158 98
rect 161 96 163 98
rect 166 96 168 98
rect 171 96 173 98
rect 176 96 178 98
rect 181 96 183 98
rect 186 96 188 98
rect 191 96 193 98
rect 196 96 198 98
rect 201 96 203 98
rect 206 96 208 98
rect 211 96 213 98
rect 216 96 218 98
rect 221 96 223 98
rect 226 96 228 98
rect 231 96 233 98
rect 236 96 238 98
rect 241 96 243 98
rect 246 96 248 98
rect 251 96 253 98
rect 256 96 258 98
rect 261 96 263 98
rect 266 96 268 98
rect 271 96 273 98
rect 276 96 278 98
rect 281 96 283 98
rect 3 93 5 95
rect 295 93 297 95
rect 3 88 5 90
rect 295 88 297 90
rect 16 86 18 88
rect 21 86 23 88
rect 26 86 28 88
rect 31 86 33 88
rect 36 86 38 88
rect 41 86 43 88
rect 46 86 48 88
rect 51 86 53 88
rect 56 86 58 88
rect 61 86 63 88
rect 66 86 68 88
rect 71 86 73 88
rect 76 86 78 88
rect 81 86 83 88
rect 86 86 88 88
rect 91 86 93 88
rect 96 86 98 88
rect 101 86 103 88
rect 106 86 108 88
rect 111 86 113 88
rect 116 86 118 88
rect 121 86 123 88
rect 126 86 128 88
rect 131 86 133 88
rect 136 86 138 88
rect 141 86 143 88
rect 146 86 148 88
rect 151 86 153 88
rect 156 86 158 88
rect 161 86 163 88
rect 166 86 168 88
rect 171 86 173 88
rect 176 86 178 88
rect 181 86 183 88
rect 186 86 188 88
rect 191 86 193 88
rect 196 86 198 88
rect 201 86 203 88
rect 206 86 208 88
rect 211 86 213 88
rect 216 86 218 88
rect 221 86 223 88
rect 226 86 228 88
rect 231 86 233 88
rect 236 86 238 88
rect 241 86 243 88
rect 246 86 248 88
rect 251 86 253 88
rect 256 86 258 88
rect 261 86 263 88
rect 266 86 268 88
rect 271 86 273 88
rect 276 86 278 88
rect 281 86 283 88
rect 3 83 5 85
rect 295 83 297 85
rect 3 78 5 80
rect 295 78 297 80
rect 16 76 18 78
rect 21 76 23 78
rect 26 76 28 78
rect 31 76 33 78
rect 36 76 38 78
rect 41 76 43 78
rect 46 76 48 78
rect 51 76 53 78
rect 56 76 58 78
rect 61 76 63 78
rect 66 76 68 78
rect 71 76 73 78
rect 76 76 78 78
rect 81 76 83 78
rect 86 76 88 78
rect 91 76 93 78
rect 96 76 98 78
rect 101 76 103 78
rect 106 76 108 78
rect 111 76 113 78
rect 116 76 118 78
rect 121 76 123 78
rect 126 76 128 78
rect 131 76 133 78
rect 136 76 138 78
rect 141 76 143 78
rect 146 76 148 78
rect 151 76 153 78
rect 156 76 158 78
rect 161 76 163 78
rect 166 76 168 78
rect 171 76 173 78
rect 176 76 178 78
rect 181 76 183 78
rect 186 76 188 78
rect 191 76 193 78
rect 196 76 198 78
rect 201 76 203 78
rect 206 76 208 78
rect 211 76 213 78
rect 216 76 218 78
rect 221 76 223 78
rect 226 76 228 78
rect 231 76 233 78
rect 236 76 238 78
rect 241 76 243 78
rect 246 76 248 78
rect 251 76 253 78
rect 256 76 258 78
rect 261 76 263 78
rect 266 76 268 78
rect 271 76 273 78
rect 276 76 278 78
rect 281 76 283 78
rect 3 73 5 75
rect 295 73 297 75
rect 3 68 5 70
rect 295 68 297 70
rect 16 66 18 68
rect 21 66 23 68
rect 26 66 28 68
rect 31 66 33 68
rect 36 66 38 68
rect 41 66 43 68
rect 46 66 48 68
rect 51 66 53 68
rect 56 66 58 68
rect 61 66 63 68
rect 66 66 68 68
rect 71 66 73 68
rect 76 66 78 68
rect 81 66 83 68
rect 86 66 88 68
rect 91 66 93 68
rect 96 66 98 68
rect 101 66 103 68
rect 106 66 108 68
rect 111 66 113 68
rect 116 66 118 68
rect 121 66 123 68
rect 126 66 128 68
rect 131 66 133 68
rect 136 66 138 68
rect 141 66 143 68
rect 146 66 148 68
rect 151 66 153 68
rect 156 66 158 68
rect 161 66 163 68
rect 166 66 168 68
rect 171 66 173 68
rect 176 66 178 68
rect 181 66 183 68
rect 186 66 188 68
rect 191 66 193 68
rect 196 66 198 68
rect 201 66 203 68
rect 206 66 208 68
rect 211 66 213 68
rect 216 66 218 68
rect 221 66 223 68
rect 226 66 228 68
rect 231 66 233 68
rect 236 66 238 68
rect 241 66 243 68
rect 246 66 248 68
rect 251 66 253 68
rect 256 66 258 68
rect 261 66 263 68
rect 266 66 268 68
rect 271 66 273 68
rect 276 66 278 68
rect 281 66 283 68
rect 3 63 5 65
rect 295 63 297 65
rect 3 58 5 60
rect 295 58 297 60
rect 16 56 18 58
rect 21 56 23 58
rect 26 56 28 58
rect 31 56 33 58
rect 36 56 38 58
rect 41 56 43 58
rect 46 56 48 58
rect 51 56 53 58
rect 56 56 58 58
rect 61 56 63 58
rect 66 56 68 58
rect 71 56 73 58
rect 76 56 78 58
rect 81 56 83 58
rect 86 56 88 58
rect 91 56 93 58
rect 96 56 98 58
rect 101 56 103 58
rect 106 56 108 58
rect 111 56 113 58
rect 116 56 118 58
rect 121 56 123 58
rect 126 56 128 58
rect 131 56 133 58
rect 136 56 138 58
rect 141 56 143 58
rect 146 56 148 58
rect 151 56 153 58
rect 156 56 158 58
rect 161 56 163 58
rect 166 56 168 58
rect 171 56 173 58
rect 176 56 178 58
rect 181 56 183 58
rect 186 56 188 58
rect 191 56 193 58
rect 196 56 198 58
rect 201 56 203 58
rect 206 56 208 58
rect 211 56 213 58
rect 216 56 218 58
rect 221 56 223 58
rect 226 56 228 58
rect 231 56 233 58
rect 236 56 238 58
rect 241 56 243 58
rect 246 56 248 58
rect 251 56 253 58
rect 256 56 258 58
rect 261 56 263 58
rect 266 56 268 58
rect 271 56 273 58
rect 276 56 278 58
rect 281 56 283 58
rect 3 53 5 55
rect 295 53 297 55
rect 3 48 5 50
rect 295 48 297 50
rect 16 46 18 48
rect 21 46 23 48
rect 26 46 28 48
rect 31 46 33 48
rect 36 46 38 48
rect 41 46 43 48
rect 46 46 48 48
rect 51 46 53 48
rect 56 46 58 48
rect 61 46 63 48
rect 66 46 68 48
rect 71 46 73 48
rect 76 46 78 48
rect 81 46 83 48
rect 86 46 88 48
rect 91 46 93 48
rect 96 46 98 48
rect 101 46 103 48
rect 106 46 108 48
rect 111 46 113 48
rect 116 46 118 48
rect 121 46 123 48
rect 126 46 128 48
rect 131 46 133 48
rect 136 46 138 48
rect 141 46 143 48
rect 146 46 148 48
rect 151 46 153 48
rect 156 46 158 48
rect 161 46 163 48
rect 166 46 168 48
rect 171 46 173 48
rect 176 46 178 48
rect 181 46 183 48
rect 186 46 188 48
rect 191 46 193 48
rect 196 46 198 48
rect 201 46 203 48
rect 206 46 208 48
rect 211 46 213 48
rect 216 46 218 48
rect 221 46 223 48
rect 226 46 228 48
rect 231 46 233 48
rect 236 46 238 48
rect 241 46 243 48
rect 246 46 248 48
rect 251 46 253 48
rect 256 46 258 48
rect 261 46 263 48
rect 266 46 268 48
rect 271 46 273 48
rect 276 46 278 48
rect 281 46 283 48
rect 3 43 5 45
rect 295 43 297 45
rect 3 38 5 40
rect 295 38 297 40
rect 16 36 18 38
rect 21 36 23 38
rect 26 36 28 38
rect 31 36 33 38
rect 36 36 38 38
rect 41 36 43 38
rect 46 36 48 38
rect 51 36 53 38
rect 56 36 58 38
rect 61 36 63 38
rect 66 36 68 38
rect 71 36 73 38
rect 76 36 78 38
rect 81 36 83 38
rect 86 36 88 38
rect 91 36 93 38
rect 96 36 98 38
rect 101 36 103 38
rect 106 36 108 38
rect 111 36 113 38
rect 116 36 118 38
rect 121 36 123 38
rect 126 36 128 38
rect 131 36 133 38
rect 136 36 138 38
rect 141 36 143 38
rect 146 36 148 38
rect 151 36 153 38
rect 156 36 158 38
rect 161 36 163 38
rect 166 36 168 38
rect 171 36 173 38
rect 176 36 178 38
rect 181 36 183 38
rect 186 36 188 38
rect 191 36 193 38
rect 196 36 198 38
rect 201 36 203 38
rect 206 36 208 38
rect 211 36 213 38
rect 216 36 218 38
rect 221 36 223 38
rect 226 36 228 38
rect 231 36 233 38
rect 236 36 238 38
rect 241 36 243 38
rect 246 36 248 38
rect 251 36 253 38
rect 256 36 258 38
rect 261 36 263 38
rect 266 36 268 38
rect 271 36 273 38
rect 276 36 278 38
rect 281 36 283 38
rect 3 33 5 35
rect 295 33 297 35
rect 3 28 5 30
rect 295 28 297 30
rect 16 26 18 28
rect 21 26 23 28
rect 26 26 28 28
rect 31 26 33 28
rect 36 26 38 28
rect 41 26 43 28
rect 46 26 48 28
rect 51 26 53 28
rect 56 26 58 28
rect 61 26 63 28
rect 66 26 68 28
rect 71 26 73 28
rect 76 26 78 28
rect 81 26 83 28
rect 86 26 88 28
rect 91 26 93 28
rect 96 26 98 28
rect 101 26 103 28
rect 106 26 108 28
rect 111 26 113 28
rect 116 26 118 28
rect 121 26 123 28
rect 126 26 128 28
rect 131 26 133 28
rect 136 26 138 28
rect 141 26 143 28
rect 146 26 148 28
rect 151 26 153 28
rect 156 26 158 28
rect 161 26 163 28
rect 166 26 168 28
rect 171 26 173 28
rect 176 26 178 28
rect 181 26 183 28
rect 186 26 188 28
rect 191 26 193 28
rect 196 26 198 28
rect 201 26 203 28
rect 206 26 208 28
rect 211 26 213 28
rect 216 26 218 28
rect 221 26 223 28
rect 226 26 228 28
rect 231 26 233 28
rect 236 26 238 28
rect 241 26 243 28
rect 246 26 248 28
rect 251 26 253 28
rect 256 26 258 28
rect 261 26 263 28
rect 266 26 268 28
rect 271 26 273 28
rect 276 26 278 28
rect 281 26 283 28
rect 3 23 5 25
rect 295 23 297 25
rect 3 18 5 20
rect 295 18 297 20
rect 16 16 18 18
rect 21 16 23 18
rect 26 16 28 18
rect 31 16 33 18
rect 36 16 38 18
rect 41 16 43 18
rect 46 16 48 18
rect 51 16 53 18
rect 56 16 58 18
rect 61 16 63 18
rect 66 16 68 18
rect 71 16 73 18
rect 76 16 78 18
rect 81 16 83 18
rect 86 16 88 18
rect 91 16 93 18
rect 96 16 98 18
rect 101 16 103 18
rect 106 16 108 18
rect 111 16 113 18
rect 116 16 118 18
rect 121 16 123 18
rect 126 16 128 18
rect 131 16 133 18
rect 136 16 138 18
rect 141 16 143 18
rect 146 16 148 18
rect 151 16 153 18
rect 156 16 158 18
rect 161 16 163 18
rect 166 16 168 18
rect 171 16 173 18
rect 176 16 178 18
rect 181 16 183 18
rect 186 16 188 18
rect 191 16 193 18
rect 196 16 198 18
rect 201 16 203 18
rect 206 16 208 18
rect 211 16 213 18
rect 216 16 218 18
rect 221 16 223 18
rect 226 16 228 18
rect 231 16 233 18
rect 236 16 238 18
rect 241 16 243 18
rect 246 16 248 18
rect 251 16 253 18
rect 256 16 258 18
rect 261 16 263 18
rect 266 16 268 18
rect 271 16 273 18
rect 276 16 278 18
rect 281 16 283 18
rect 3 13 5 15
rect 295 13 297 15
rect 3 8 5 10
rect 295 8 297 10
rect 3 3 5 5
rect 11 3 13 5
rect 16 3 18 5
rect 21 3 23 5
rect 26 3 28 5
rect 31 3 33 5
rect 36 3 38 5
rect 41 3 43 5
rect 46 3 48 5
rect 51 3 53 5
rect 56 3 58 5
rect 61 3 63 5
rect 66 3 68 5
rect 71 3 73 5
rect 76 3 78 5
rect 81 3 83 5
rect 86 3 88 5
rect 91 3 93 5
rect 207 3 209 5
rect 212 3 214 5
rect 217 3 219 5
rect 222 3 224 5
rect 227 3 229 5
rect 232 3 234 5
rect 237 3 239 5
rect 242 3 244 5
rect 247 3 249 5
rect 252 3 254 5
rect 257 3 259 5
rect 262 3 264 5
rect 267 3 269 5
rect 272 3 274 5
rect 277 3 279 5
rect 282 3 284 5
rect 287 3 289 5
rect 295 3 297 5
<< metal1 >>
rect 20 740 280 1000
rect 62 730 238 740
rect 72 720 228 730
rect 82 710 218 720
rect 92 700 208 710
rect 102 670 198 700
rect 0 659 300 670
rect 0 423 11 659
rect 102 653 198 659
rect 36 649 120 650
rect 20 621 120 649
rect 20 590 51 621
rect 123 618 177 653
rect 180 621 280 650
rect 56 593 140 618
rect 20 557 120 590
rect 123 588 140 593
rect 143 591 157 615
rect 160 593 244 618
rect 160 588 177 593
rect 249 590 280 621
rect 20 526 51 557
rect 123 554 177 588
rect 180 557 280 590
rect 56 529 140 554
rect 20 492 120 526
rect 123 524 140 529
rect 143 527 157 551
rect 160 529 244 554
rect 160 524 177 529
rect 249 526 280 557
rect 20 461 51 492
rect 123 489 177 524
rect 180 492 280 526
rect 56 464 140 489
rect 20 432 120 461
rect 123 459 140 464
rect 143 462 157 486
rect 160 464 244 489
rect 160 459 177 464
rect 249 461 280 492
rect 123 429 177 459
rect 180 432 280 461
rect 102 423 198 429
rect 289 423 300 659
rect 0 344 300 423
rect 102 329 198 344
rect 0 252 99 326
rect 0 7 7 252
rect 102 246 140 329
rect 143 252 157 326
rect 160 246 198 329
rect 201 252 300 326
rect 102 245 198 246
rect 15 15 285 245
rect 0 1 99 7
rect 102 -11 198 15
rect 293 7 300 252
rect 201 1 300 7
<< metal2 >>
rect 20 740 280 1000
rect 0 440 300 670
rect 0 344 300 424
rect 0 246 300 326
rect 0 0 300 230
<< gv1 >>
rect 41 977 43 979
rect 53 977 55 979
rect 65 977 67 979
rect 77 977 79 979
rect 89 977 91 979
rect 101 977 103 979
rect 113 977 115 979
rect 125 977 127 979
rect 137 977 139 979
rect 149 977 151 979
rect 161 977 163 979
rect 173 977 175 979
rect 185 977 187 979
rect 197 977 199 979
rect 209 977 211 979
rect 221 977 223 979
rect 233 977 235 979
rect 245 977 247 979
rect 257 977 259 979
rect 41 965 43 967
rect 53 965 55 967
rect 65 965 67 967
rect 77 965 79 967
rect 89 965 91 967
rect 101 965 103 967
rect 113 965 115 967
rect 125 965 127 967
rect 137 965 139 967
rect 149 965 151 967
rect 161 965 163 967
rect 173 965 175 967
rect 185 965 187 967
rect 197 965 199 967
rect 209 965 211 967
rect 221 965 223 967
rect 233 965 235 967
rect 245 965 247 967
rect 257 965 259 967
rect 41 953 43 955
rect 53 953 55 955
rect 65 953 67 955
rect 77 953 79 955
rect 89 953 91 955
rect 101 953 103 955
rect 113 953 115 955
rect 125 953 127 955
rect 137 953 139 955
rect 149 953 151 955
rect 161 953 163 955
rect 173 953 175 955
rect 185 953 187 955
rect 197 953 199 955
rect 209 953 211 955
rect 221 953 223 955
rect 233 953 235 955
rect 245 953 247 955
rect 257 953 259 955
rect 41 941 43 943
rect 53 941 55 943
rect 65 941 67 943
rect 77 941 79 943
rect 89 941 91 943
rect 101 941 103 943
rect 113 941 115 943
rect 125 941 127 943
rect 137 941 139 943
rect 149 941 151 943
rect 161 941 163 943
rect 173 941 175 943
rect 185 941 187 943
rect 197 941 199 943
rect 209 941 211 943
rect 221 941 223 943
rect 233 941 235 943
rect 245 941 247 943
rect 257 941 259 943
rect 41 929 43 931
rect 53 929 55 931
rect 65 929 67 931
rect 77 929 79 931
rect 89 929 91 931
rect 101 929 103 931
rect 113 929 115 931
rect 125 929 127 931
rect 137 929 139 931
rect 149 929 151 931
rect 161 929 163 931
rect 173 929 175 931
rect 185 929 187 931
rect 197 929 199 931
rect 209 929 211 931
rect 221 929 223 931
rect 233 929 235 931
rect 245 929 247 931
rect 257 929 259 931
rect 41 917 43 919
rect 53 917 55 919
rect 65 917 67 919
rect 77 917 79 919
rect 89 917 91 919
rect 101 917 103 919
rect 113 917 115 919
rect 125 917 127 919
rect 137 917 139 919
rect 149 917 151 919
rect 161 917 163 919
rect 173 917 175 919
rect 185 917 187 919
rect 197 917 199 919
rect 209 917 211 919
rect 221 917 223 919
rect 233 917 235 919
rect 245 917 247 919
rect 257 917 259 919
rect 41 905 43 907
rect 53 905 55 907
rect 65 905 67 907
rect 77 905 79 907
rect 89 905 91 907
rect 101 905 103 907
rect 113 905 115 907
rect 125 905 127 907
rect 137 905 139 907
rect 149 905 151 907
rect 161 905 163 907
rect 173 905 175 907
rect 185 905 187 907
rect 197 905 199 907
rect 209 905 211 907
rect 221 905 223 907
rect 233 905 235 907
rect 245 905 247 907
rect 257 905 259 907
rect 41 893 43 895
rect 53 893 55 895
rect 65 893 67 895
rect 77 893 79 895
rect 89 893 91 895
rect 101 893 103 895
rect 113 893 115 895
rect 125 893 127 895
rect 137 893 139 895
rect 149 893 151 895
rect 161 893 163 895
rect 173 893 175 895
rect 185 893 187 895
rect 197 893 199 895
rect 209 893 211 895
rect 221 893 223 895
rect 233 893 235 895
rect 245 893 247 895
rect 257 893 259 895
rect 41 881 43 883
rect 53 881 55 883
rect 65 881 67 883
rect 77 881 79 883
rect 89 881 91 883
rect 101 881 103 883
rect 113 881 115 883
rect 125 881 127 883
rect 137 881 139 883
rect 149 881 151 883
rect 161 881 163 883
rect 173 881 175 883
rect 185 881 187 883
rect 197 881 199 883
rect 209 881 211 883
rect 221 881 223 883
rect 233 881 235 883
rect 245 881 247 883
rect 257 881 259 883
rect 41 869 43 871
rect 53 869 55 871
rect 65 869 67 871
rect 77 869 79 871
rect 89 869 91 871
rect 101 869 103 871
rect 113 869 115 871
rect 125 869 127 871
rect 137 869 139 871
rect 149 869 151 871
rect 161 869 163 871
rect 173 869 175 871
rect 185 869 187 871
rect 197 869 199 871
rect 209 869 211 871
rect 221 869 223 871
rect 233 869 235 871
rect 245 869 247 871
rect 257 869 259 871
rect 41 857 43 859
rect 53 857 55 859
rect 65 857 67 859
rect 77 857 79 859
rect 89 857 91 859
rect 101 857 103 859
rect 113 857 115 859
rect 125 857 127 859
rect 137 857 139 859
rect 149 857 151 859
rect 161 857 163 859
rect 173 857 175 859
rect 185 857 187 859
rect 197 857 199 859
rect 209 857 211 859
rect 221 857 223 859
rect 233 857 235 859
rect 245 857 247 859
rect 257 857 259 859
rect 41 845 43 847
rect 53 845 55 847
rect 65 845 67 847
rect 77 845 79 847
rect 89 845 91 847
rect 101 845 103 847
rect 113 845 115 847
rect 125 845 127 847
rect 137 845 139 847
rect 149 845 151 847
rect 161 845 163 847
rect 173 845 175 847
rect 185 845 187 847
rect 197 845 199 847
rect 209 845 211 847
rect 221 845 223 847
rect 233 845 235 847
rect 245 845 247 847
rect 257 845 259 847
rect 41 833 43 835
rect 53 833 55 835
rect 65 833 67 835
rect 77 833 79 835
rect 89 833 91 835
rect 101 833 103 835
rect 113 833 115 835
rect 125 833 127 835
rect 137 833 139 835
rect 149 833 151 835
rect 161 833 163 835
rect 173 833 175 835
rect 185 833 187 835
rect 197 833 199 835
rect 209 833 211 835
rect 221 833 223 835
rect 233 833 235 835
rect 245 833 247 835
rect 257 833 259 835
rect 41 821 43 823
rect 53 821 55 823
rect 65 821 67 823
rect 77 821 79 823
rect 89 821 91 823
rect 101 821 103 823
rect 113 821 115 823
rect 125 821 127 823
rect 137 821 139 823
rect 149 821 151 823
rect 161 821 163 823
rect 173 821 175 823
rect 185 821 187 823
rect 197 821 199 823
rect 209 821 211 823
rect 221 821 223 823
rect 233 821 235 823
rect 245 821 247 823
rect 257 821 259 823
rect 41 809 43 811
rect 53 809 55 811
rect 65 809 67 811
rect 77 809 79 811
rect 89 809 91 811
rect 101 809 103 811
rect 113 809 115 811
rect 125 809 127 811
rect 137 809 139 811
rect 149 809 151 811
rect 161 809 163 811
rect 173 809 175 811
rect 185 809 187 811
rect 197 809 199 811
rect 209 809 211 811
rect 221 809 223 811
rect 233 809 235 811
rect 245 809 247 811
rect 257 809 259 811
rect 41 797 43 799
rect 53 797 55 799
rect 65 797 67 799
rect 77 797 79 799
rect 89 797 91 799
rect 101 797 103 799
rect 113 797 115 799
rect 125 797 127 799
rect 137 797 139 799
rect 149 797 151 799
rect 161 797 163 799
rect 173 797 175 799
rect 185 797 187 799
rect 197 797 199 799
rect 209 797 211 799
rect 221 797 223 799
rect 233 797 235 799
rect 245 797 247 799
rect 257 797 259 799
rect 41 785 43 787
rect 53 785 55 787
rect 65 785 67 787
rect 77 785 79 787
rect 89 785 91 787
rect 101 785 103 787
rect 113 785 115 787
rect 125 785 127 787
rect 137 785 139 787
rect 149 785 151 787
rect 161 785 163 787
rect 173 785 175 787
rect 185 785 187 787
rect 197 785 199 787
rect 209 785 211 787
rect 221 785 223 787
rect 233 785 235 787
rect 245 785 247 787
rect 257 785 259 787
rect 41 773 43 775
rect 53 773 55 775
rect 65 773 67 775
rect 77 773 79 775
rect 89 773 91 775
rect 101 773 103 775
rect 113 773 115 775
rect 125 773 127 775
rect 137 773 139 775
rect 149 773 151 775
rect 161 773 163 775
rect 173 773 175 775
rect 185 773 187 775
rect 197 773 199 775
rect 209 773 211 775
rect 221 773 223 775
rect 233 773 235 775
rect 245 773 247 775
rect 257 773 259 775
rect 41 761 43 763
rect 53 761 55 763
rect 65 761 67 763
rect 77 761 79 763
rect 89 761 91 763
rect 101 761 103 763
rect 113 761 115 763
rect 125 761 127 763
rect 137 761 139 763
rect 149 761 151 763
rect 161 761 163 763
rect 173 761 175 763
rect 185 761 187 763
rect 197 761 199 763
rect 209 761 211 763
rect 221 761 223 763
rect 233 761 235 763
rect 245 761 247 763
rect 257 761 259 763
rect 22 646 24 648
rect 276 646 278 648
rect 22 641 24 643
rect 276 641 278 643
rect 37 639 39 641
rect 42 639 44 641
rect 47 639 49 641
rect 52 639 54 641
rect 57 639 59 641
rect 62 639 64 641
rect 67 639 69 641
rect 72 639 74 641
rect 77 639 79 641
rect 82 639 84 641
rect 87 639 89 641
rect 92 639 94 641
rect 97 639 99 641
rect 102 639 104 641
rect 107 639 109 641
rect 112 639 114 641
rect 117 639 119 641
rect 181 639 183 641
rect 186 639 188 641
rect 191 639 193 641
rect 196 639 198 641
rect 201 639 203 641
rect 206 639 208 641
rect 211 639 213 641
rect 216 639 218 641
rect 221 639 223 641
rect 226 639 228 641
rect 231 639 233 641
rect 236 639 238 641
rect 241 639 243 641
rect 246 639 248 641
rect 251 639 253 641
rect 256 639 258 641
rect 261 639 263 641
rect 22 636 24 638
rect 276 636 278 638
rect 22 631 24 633
rect 276 631 278 633
rect 22 626 24 628
rect 276 626 278 628
rect 22 621 24 623
rect 40 622 42 624
rect 45 622 47 624
rect 53 622 55 624
rect 58 622 60 624
rect 63 622 65 624
rect 68 622 70 624
rect 73 622 75 624
rect 78 622 80 624
rect 83 622 85 624
rect 88 622 90 624
rect 93 622 95 624
rect 98 622 100 624
rect 103 622 105 624
rect 108 622 110 624
rect 113 622 115 624
rect 185 622 187 624
rect 190 622 192 624
rect 195 622 197 624
rect 200 622 202 624
rect 205 622 207 624
rect 210 622 212 624
rect 215 622 217 624
rect 220 622 222 624
rect 225 622 227 624
rect 230 622 232 624
rect 235 622 237 624
rect 240 622 242 624
rect 245 622 247 624
rect 253 622 255 624
rect 258 622 260 624
rect 276 621 278 623
rect 22 616 24 618
rect 40 617 42 619
rect 45 617 47 619
rect 253 617 255 619
rect 258 617 260 619
rect 276 616 278 618
rect 22 611 24 613
rect 40 612 42 614
rect 45 612 47 614
rect 253 612 255 614
rect 258 612 260 614
rect 276 611 278 613
rect 22 606 24 608
rect 40 607 42 609
rect 45 607 47 609
rect 144 607 146 609
rect 149 607 151 609
rect 154 607 156 609
rect 253 607 255 609
rect 258 607 260 609
rect 276 606 278 608
rect 22 601 24 603
rect 40 602 42 604
rect 45 602 47 604
rect 253 602 255 604
rect 258 602 260 604
rect 276 601 278 603
rect 22 596 24 598
rect 40 597 42 599
rect 45 597 47 599
rect 144 597 146 599
rect 149 597 151 599
rect 154 597 156 599
rect 253 597 255 599
rect 258 597 260 599
rect 276 596 278 598
rect 22 591 24 593
rect 40 592 42 594
rect 45 592 47 594
rect 253 592 255 594
rect 258 592 260 594
rect 276 591 278 593
rect 22 586 24 588
rect 40 587 42 589
rect 45 587 47 589
rect 53 587 55 589
rect 58 587 60 589
rect 63 587 65 589
rect 68 587 70 589
rect 73 587 75 589
rect 78 587 80 589
rect 83 587 85 589
rect 88 587 90 589
rect 93 587 95 589
rect 98 587 100 589
rect 103 587 105 589
rect 108 587 110 589
rect 113 587 115 589
rect 185 587 187 589
rect 190 587 192 589
rect 195 587 197 589
rect 200 587 202 589
rect 205 587 207 589
rect 210 587 212 589
rect 215 587 217 589
rect 220 587 222 589
rect 225 587 227 589
rect 230 587 232 589
rect 235 587 237 589
rect 240 587 242 589
rect 245 587 247 589
rect 253 587 255 589
rect 258 587 260 589
rect 276 586 278 588
rect 22 581 24 583
rect 276 581 278 583
rect 22 576 24 578
rect 276 576 278 578
rect 22 571 24 573
rect 276 571 278 573
rect 22 566 24 568
rect 276 566 278 568
rect 22 561 24 563
rect 276 561 278 563
rect 40 558 42 560
rect 45 558 47 560
rect 53 558 55 560
rect 58 558 60 560
rect 63 558 65 560
rect 68 558 70 560
rect 73 558 75 560
rect 78 558 80 560
rect 83 558 85 560
rect 88 558 90 560
rect 93 558 95 560
rect 98 558 100 560
rect 103 558 105 560
rect 108 558 110 560
rect 113 558 115 560
rect 185 558 187 560
rect 190 558 192 560
rect 195 558 197 560
rect 200 558 202 560
rect 205 558 207 560
rect 210 558 212 560
rect 215 558 217 560
rect 220 558 222 560
rect 225 558 227 560
rect 230 558 232 560
rect 235 558 237 560
rect 240 558 242 560
rect 245 558 247 560
rect 253 558 255 560
rect 258 558 260 560
rect 22 556 24 558
rect 276 556 278 558
rect 40 553 42 555
rect 45 553 47 555
rect 253 553 255 555
rect 258 553 260 555
rect 22 551 24 553
rect 276 551 278 553
rect 40 548 42 550
rect 45 548 47 550
rect 253 548 255 550
rect 258 548 260 550
rect 22 546 24 548
rect 276 546 278 548
rect 40 543 42 545
rect 45 543 47 545
rect 144 543 146 545
rect 149 543 151 545
rect 154 543 156 545
rect 253 543 255 545
rect 258 543 260 545
rect 22 541 24 543
rect 276 541 278 543
rect 40 538 42 540
rect 45 538 47 540
rect 253 538 255 540
rect 258 538 260 540
rect 22 536 24 538
rect 276 536 278 538
rect 40 533 42 535
rect 45 533 47 535
rect 144 533 146 535
rect 149 533 151 535
rect 154 533 156 535
rect 253 533 255 535
rect 258 533 260 535
rect 22 531 24 533
rect 276 531 278 533
rect 40 528 42 530
rect 45 528 47 530
rect 253 528 255 530
rect 258 528 260 530
rect 22 526 24 528
rect 276 526 278 528
rect 40 523 42 525
rect 45 523 47 525
rect 53 523 55 525
rect 58 523 60 525
rect 63 523 65 525
rect 68 523 70 525
rect 73 523 75 525
rect 78 523 80 525
rect 83 523 85 525
rect 88 523 90 525
rect 93 523 95 525
rect 98 523 100 525
rect 103 523 105 525
rect 108 523 110 525
rect 113 523 115 525
rect 185 523 187 525
rect 190 523 192 525
rect 195 523 197 525
rect 200 523 202 525
rect 205 523 207 525
rect 210 523 212 525
rect 215 523 217 525
rect 220 523 222 525
rect 225 523 227 525
rect 230 523 232 525
rect 235 523 237 525
rect 240 523 242 525
rect 245 523 247 525
rect 253 523 255 525
rect 258 523 260 525
rect 22 521 24 523
rect 276 521 278 523
rect 22 516 24 518
rect 276 516 278 518
rect 22 511 24 513
rect 276 511 278 513
rect 22 506 24 508
rect 276 506 278 508
rect 22 501 24 503
rect 276 501 278 503
rect 22 496 24 498
rect 276 496 278 498
rect 40 493 42 495
rect 45 493 47 495
rect 53 493 55 495
rect 58 493 60 495
rect 63 493 65 495
rect 68 493 70 495
rect 73 493 75 495
rect 78 493 80 495
rect 83 493 85 495
rect 88 493 90 495
rect 93 493 95 495
rect 98 493 100 495
rect 103 493 105 495
rect 108 493 110 495
rect 113 493 115 495
rect 185 493 187 495
rect 190 493 192 495
rect 195 493 197 495
rect 200 493 202 495
rect 205 493 207 495
rect 210 493 212 495
rect 215 493 217 495
rect 220 493 222 495
rect 225 493 227 495
rect 230 493 232 495
rect 235 493 237 495
rect 240 493 242 495
rect 245 493 247 495
rect 253 493 255 495
rect 258 493 260 495
rect 22 491 24 493
rect 276 491 278 493
rect 40 488 42 490
rect 45 488 47 490
rect 253 488 255 490
rect 258 488 260 490
rect 22 486 24 488
rect 276 486 278 488
rect 40 483 42 485
rect 45 483 47 485
rect 253 483 255 485
rect 258 483 260 485
rect 22 481 24 483
rect 276 481 278 483
rect 40 478 42 480
rect 45 478 47 480
rect 144 478 146 480
rect 149 478 151 480
rect 154 478 156 480
rect 253 478 255 480
rect 258 478 260 480
rect 22 476 24 478
rect 276 476 278 478
rect 40 473 42 475
rect 45 473 47 475
rect 253 473 255 475
rect 258 473 260 475
rect 22 471 24 473
rect 276 471 278 473
rect 40 468 42 470
rect 45 468 47 470
rect 144 468 146 470
rect 149 468 151 470
rect 154 468 156 470
rect 253 468 255 470
rect 258 468 260 470
rect 22 466 24 468
rect 276 466 278 468
rect 40 463 42 465
rect 45 463 47 465
rect 253 463 255 465
rect 258 463 260 465
rect 22 461 24 463
rect 276 461 278 463
rect 40 458 42 460
rect 45 458 47 460
rect 53 458 55 460
rect 58 458 60 460
rect 63 458 65 460
rect 68 458 70 460
rect 73 458 75 460
rect 78 458 80 460
rect 83 458 85 460
rect 88 458 90 460
rect 93 458 95 460
rect 98 458 100 460
rect 103 458 105 460
rect 108 458 110 460
rect 113 458 115 460
rect 185 458 187 460
rect 190 458 192 460
rect 195 458 197 460
rect 200 458 202 460
rect 205 458 207 460
rect 210 458 212 460
rect 215 458 217 460
rect 220 458 222 460
rect 225 458 227 460
rect 230 458 232 460
rect 235 458 237 460
rect 240 458 242 460
rect 245 458 247 460
rect 253 458 255 460
rect 258 458 260 460
rect 22 456 24 458
rect 276 456 278 458
rect 22 451 24 453
rect 276 451 278 453
rect 22 446 24 448
rect 276 446 278 448
rect 4 410 6 412
rect 9 410 11 412
rect 14 410 16 412
rect 19 410 21 412
rect 24 410 26 412
rect 29 410 31 412
rect 34 410 36 412
rect 39 410 41 412
rect 44 410 46 412
rect 49 410 51 412
rect 54 410 56 412
rect 59 410 61 412
rect 64 410 66 412
rect 69 410 71 412
rect 74 410 76 412
rect 79 410 81 412
rect 84 410 86 412
rect 89 410 91 412
rect 94 410 96 412
rect 99 410 101 412
rect 104 410 106 412
rect 109 410 111 412
rect 114 410 116 412
rect 119 410 121 412
rect 124 410 126 412
rect 129 410 131 412
rect 134 410 136 412
rect 139 410 141 412
rect 144 410 146 412
rect 149 410 151 412
rect 154 410 156 412
rect 159 410 161 412
rect 164 410 166 412
rect 169 410 171 412
rect 174 410 176 412
rect 179 410 181 412
rect 184 410 186 412
rect 189 410 191 412
rect 194 410 196 412
rect 199 410 201 412
rect 204 410 206 412
rect 209 410 211 412
rect 214 410 216 412
rect 219 410 221 412
rect 224 410 226 412
rect 229 410 231 412
rect 234 410 236 412
rect 239 410 241 412
rect 244 410 246 412
rect 249 410 251 412
rect 254 410 256 412
rect 259 410 261 412
rect 264 410 266 412
rect 269 410 271 412
rect 274 410 276 412
rect 279 410 281 412
rect 284 410 286 412
rect 289 410 291 412
rect 294 410 296 412
rect 4 400 6 402
rect 9 400 11 402
rect 14 400 16 402
rect 19 400 21 402
rect 24 400 26 402
rect 29 400 31 402
rect 34 400 36 402
rect 39 400 41 402
rect 44 400 46 402
rect 49 400 51 402
rect 54 400 56 402
rect 59 400 61 402
rect 64 400 66 402
rect 69 400 71 402
rect 74 400 76 402
rect 79 400 81 402
rect 84 400 86 402
rect 89 400 91 402
rect 94 400 96 402
rect 99 400 101 402
rect 104 400 106 402
rect 109 400 111 402
rect 114 400 116 402
rect 119 400 121 402
rect 124 400 126 402
rect 129 400 131 402
rect 134 400 136 402
rect 139 400 141 402
rect 144 400 146 402
rect 149 400 151 402
rect 154 400 156 402
rect 159 400 161 402
rect 164 400 166 402
rect 169 400 171 402
rect 174 400 176 402
rect 179 400 181 402
rect 184 400 186 402
rect 189 400 191 402
rect 194 400 196 402
rect 199 400 201 402
rect 204 400 206 402
rect 209 400 211 402
rect 214 400 216 402
rect 219 400 221 402
rect 224 400 226 402
rect 229 400 231 402
rect 234 400 236 402
rect 239 400 241 402
rect 244 400 246 402
rect 249 400 251 402
rect 254 400 256 402
rect 259 400 261 402
rect 264 400 266 402
rect 269 400 271 402
rect 274 400 276 402
rect 279 400 281 402
rect 284 400 286 402
rect 289 400 291 402
rect 294 400 296 402
rect 4 390 6 392
rect 9 390 11 392
rect 14 390 16 392
rect 19 390 21 392
rect 24 390 26 392
rect 29 390 31 392
rect 34 390 36 392
rect 39 390 41 392
rect 44 390 46 392
rect 49 390 51 392
rect 54 390 56 392
rect 59 390 61 392
rect 64 390 66 392
rect 69 390 71 392
rect 74 390 76 392
rect 79 390 81 392
rect 84 390 86 392
rect 89 390 91 392
rect 94 390 96 392
rect 99 390 101 392
rect 104 390 106 392
rect 109 390 111 392
rect 114 390 116 392
rect 119 390 121 392
rect 124 390 126 392
rect 129 390 131 392
rect 134 390 136 392
rect 139 390 141 392
rect 144 390 146 392
rect 149 390 151 392
rect 154 390 156 392
rect 159 390 161 392
rect 164 390 166 392
rect 169 390 171 392
rect 174 390 176 392
rect 179 390 181 392
rect 184 390 186 392
rect 189 390 191 392
rect 194 390 196 392
rect 199 390 201 392
rect 204 390 206 392
rect 209 390 211 392
rect 214 390 216 392
rect 219 390 221 392
rect 224 390 226 392
rect 229 390 231 392
rect 234 390 236 392
rect 239 390 241 392
rect 244 390 246 392
rect 249 390 251 392
rect 254 390 256 392
rect 259 390 261 392
rect 264 390 266 392
rect 269 390 271 392
rect 274 390 276 392
rect 279 390 281 392
rect 284 390 286 392
rect 289 390 291 392
rect 294 390 296 392
rect 4 380 6 382
rect 9 380 11 382
rect 14 380 16 382
rect 19 380 21 382
rect 24 380 26 382
rect 29 380 31 382
rect 34 380 36 382
rect 39 380 41 382
rect 44 380 46 382
rect 49 380 51 382
rect 54 380 56 382
rect 59 380 61 382
rect 64 380 66 382
rect 69 380 71 382
rect 74 380 76 382
rect 79 380 81 382
rect 84 380 86 382
rect 89 380 91 382
rect 94 380 96 382
rect 99 380 101 382
rect 104 380 106 382
rect 109 380 111 382
rect 114 380 116 382
rect 119 380 121 382
rect 124 380 126 382
rect 129 380 131 382
rect 134 380 136 382
rect 139 380 141 382
rect 144 380 146 382
rect 149 380 151 382
rect 154 380 156 382
rect 159 380 161 382
rect 164 380 166 382
rect 169 380 171 382
rect 174 380 176 382
rect 179 380 181 382
rect 184 380 186 382
rect 189 380 191 382
rect 194 380 196 382
rect 199 380 201 382
rect 204 380 206 382
rect 209 380 211 382
rect 214 380 216 382
rect 219 380 221 382
rect 224 380 226 382
rect 229 380 231 382
rect 234 380 236 382
rect 239 380 241 382
rect 244 380 246 382
rect 249 380 251 382
rect 254 380 256 382
rect 259 380 261 382
rect 264 380 266 382
rect 269 380 271 382
rect 274 380 276 382
rect 279 380 281 382
rect 284 380 286 382
rect 289 380 291 382
rect 294 380 296 382
rect 4 370 6 372
rect 9 370 11 372
rect 14 370 16 372
rect 19 370 21 372
rect 24 370 26 372
rect 29 370 31 372
rect 34 370 36 372
rect 39 370 41 372
rect 44 370 46 372
rect 49 370 51 372
rect 54 370 56 372
rect 59 370 61 372
rect 64 370 66 372
rect 69 370 71 372
rect 74 370 76 372
rect 79 370 81 372
rect 84 370 86 372
rect 89 370 91 372
rect 94 370 96 372
rect 99 370 101 372
rect 104 370 106 372
rect 109 370 111 372
rect 114 370 116 372
rect 119 370 121 372
rect 124 370 126 372
rect 129 370 131 372
rect 134 370 136 372
rect 139 370 141 372
rect 144 370 146 372
rect 149 370 151 372
rect 154 370 156 372
rect 159 370 161 372
rect 164 370 166 372
rect 169 370 171 372
rect 174 370 176 372
rect 179 370 181 372
rect 184 370 186 372
rect 189 370 191 372
rect 194 370 196 372
rect 199 370 201 372
rect 204 370 206 372
rect 209 370 211 372
rect 214 370 216 372
rect 219 370 221 372
rect 224 370 226 372
rect 229 370 231 372
rect 234 370 236 372
rect 239 370 241 372
rect 244 370 246 372
rect 249 370 251 372
rect 254 370 256 372
rect 259 370 261 372
rect 264 370 266 372
rect 269 370 271 372
rect 274 370 276 372
rect 279 370 281 372
rect 284 370 286 372
rect 289 370 291 372
rect 294 370 296 372
rect 4 360 6 362
rect 9 360 11 362
rect 14 360 16 362
rect 19 360 21 362
rect 24 360 26 362
rect 29 360 31 362
rect 34 360 36 362
rect 39 360 41 362
rect 44 360 46 362
rect 49 360 51 362
rect 54 360 56 362
rect 59 360 61 362
rect 64 360 66 362
rect 69 360 71 362
rect 74 360 76 362
rect 79 360 81 362
rect 84 360 86 362
rect 89 360 91 362
rect 94 360 96 362
rect 99 360 101 362
rect 104 360 106 362
rect 109 360 111 362
rect 114 360 116 362
rect 119 360 121 362
rect 124 360 126 362
rect 129 360 131 362
rect 134 360 136 362
rect 139 360 141 362
rect 144 360 146 362
rect 149 360 151 362
rect 154 360 156 362
rect 159 360 161 362
rect 164 360 166 362
rect 169 360 171 362
rect 174 360 176 362
rect 179 360 181 362
rect 184 360 186 362
rect 189 360 191 362
rect 194 360 196 362
rect 199 360 201 362
rect 204 360 206 362
rect 209 360 211 362
rect 214 360 216 362
rect 219 360 221 362
rect 224 360 226 362
rect 229 360 231 362
rect 234 360 236 362
rect 239 360 241 362
rect 244 360 246 362
rect 249 360 251 362
rect 254 360 256 362
rect 259 360 261 362
rect 264 360 266 362
rect 269 360 271 362
rect 274 360 276 362
rect 279 360 281 362
rect 284 360 286 362
rect 289 360 291 362
rect 294 360 296 362
rect 4 350 6 352
rect 9 350 11 352
rect 14 350 16 352
rect 19 350 21 352
rect 24 350 26 352
rect 29 350 31 352
rect 34 350 36 352
rect 39 350 41 352
rect 44 350 46 352
rect 49 350 51 352
rect 54 350 56 352
rect 59 350 61 352
rect 64 350 66 352
rect 69 350 71 352
rect 74 350 76 352
rect 79 350 81 352
rect 84 350 86 352
rect 89 350 91 352
rect 94 350 96 352
rect 99 350 101 352
rect 104 350 106 352
rect 109 350 111 352
rect 114 350 116 352
rect 119 350 121 352
rect 124 350 126 352
rect 129 350 131 352
rect 134 350 136 352
rect 139 350 141 352
rect 144 350 146 352
rect 149 350 151 352
rect 154 350 156 352
rect 159 350 161 352
rect 164 350 166 352
rect 169 350 171 352
rect 174 350 176 352
rect 179 350 181 352
rect 184 350 186 352
rect 189 350 191 352
rect 194 350 196 352
rect 199 350 201 352
rect 204 350 206 352
rect 209 350 211 352
rect 214 350 216 352
rect 219 350 221 352
rect 224 350 226 352
rect 229 350 231 352
rect 234 350 236 352
rect 239 350 241 352
rect 244 350 246 352
rect 249 350 251 352
rect 254 350 256 352
rect 259 350 261 352
rect 264 350 266 352
rect 269 350 271 352
rect 274 350 276 352
rect 279 350 281 352
rect 284 350 286 352
rect 289 350 291 352
rect 294 350 296 352
rect 3 318 5 320
rect 8 318 10 320
rect 13 318 15 320
rect 18 318 20 320
rect 23 318 25 320
rect 28 318 30 320
rect 33 318 35 320
rect 38 318 40 320
rect 43 318 45 320
rect 48 318 50 320
rect 53 318 55 320
rect 58 318 60 320
rect 63 318 65 320
rect 68 318 70 320
rect 73 318 75 320
rect 78 318 80 320
rect 83 318 85 320
rect 88 318 90 320
rect 93 318 95 320
rect 144 318 146 320
rect 149 318 151 320
rect 154 318 156 320
rect 205 318 207 320
rect 210 318 212 320
rect 215 318 217 320
rect 220 318 222 320
rect 225 318 227 320
rect 230 318 232 320
rect 235 318 237 320
rect 240 318 242 320
rect 245 318 247 320
rect 250 318 252 320
rect 255 318 257 320
rect 260 318 262 320
rect 265 318 267 320
rect 270 318 272 320
rect 275 318 277 320
rect 280 318 282 320
rect 285 318 287 320
rect 290 318 292 320
rect 295 318 297 320
rect 3 308 5 310
rect 8 308 10 310
rect 13 308 15 310
rect 18 308 20 310
rect 23 308 25 310
rect 28 308 30 310
rect 33 308 35 310
rect 38 308 40 310
rect 43 308 45 310
rect 48 308 50 310
rect 53 308 55 310
rect 58 308 60 310
rect 63 308 65 310
rect 68 308 70 310
rect 73 308 75 310
rect 78 308 80 310
rect 83 308 85 310
rect 88 308 90 310
rect 93 308 95 310
rect 144 308 146 310
rect 149 308 151 310
rect 154 308 156 310
rect 205 308 207 310
rect 210 308 212 310
rect 215 308 217 310
rect 220 308 222 310
rect 225 308 227 310
rect 230 308 232 310
rect 235 308 237 310
rect 240 308 242 310
rect 245 308 247 310
rect 250 308 252 310
rect 255 308 257 310
rect 260 308 262 310
rect 265 308 267 310
rect 270 308 272 310
rect 275 308 277 310
rect 280 308 282 310
rect 285 308 287 310
rect 290 308 292 310
rect 295 308 297 310
rect 3 298 5 300
rect 8 298 10 300
rect 13 298 15 300
rect 18 298 20 300
rect 23 298 25 300
rect 28 298 30 300
rect 33 298 35 300
rect 38 298 40 300
rect 43 298 45 300
rect 48 298 50 300
rect 53 298 55 300
rect 58 298 60 300
rect 63 298 65 300
rect 68 298 70 300
rect 73 298 75 300
rect 78 298 80 300
rect 83 298 85 300
rect 88 298 90 300
rect 93 298 95 300
rect 144 298 146 300
rect 149 298 151 300
rect 154 298 156 300
rect 205 298 207 300
rect 210 298 212 300
rect 215 298 217 300
rect 220 298 222 300
rect 225 298 227 300
rect 230 298 232 300
rect 235 298 237 300
rect 240 298 242 300
rect 245 298 247 300
rect 250 298 252 300
rect 255 298 257 300
rect 260 298 262 300
rect 265 298 267 300
rect 270 298 272 300
rect 275 298 277 300
rect 280 298 282 300
rect 285 298 287 300
rect 290 298 292 300
rect 295 298 297 300
rect 3 288 5 290
rect 8 288 10 290
rect 13 288 15 290
rect 18 288 20 290
rect 23 288 25 290
rect 28 288 30 290
rect 33 288 35 290
rect 38 288 40 290
rect 43 288 45 290
rect 48 288 50 290
rect 53 288 55 290
rect 58 288 60 290
rect 63 288 65 290
rect 68 288 70 290
rect 73 288 75 290
rect 78 288 80 290
rect 83 288 85 290
rect 88 288 90 290
rect 93 288 95 290
rect 144 288 146 290
rect 149 288 151 290
rect 154 288 156 290
rect 205 288 207 290
rect 210 288 212 290
rect 215 288 217 290
rect 220 288 222 290
rect 225 288 227 290
rect 230 288 232 290
rect 235 288 237 290
rect 240 288 242 290
rect 245 288 247 290
rect 250 288 252 290
rect 255 288 257 290
rect 260 288 262 290
rect 265 288 267 290
rect 270 288 272 290
rect 275 288 277 290
rect 280 288 282 290
rect 285 288 287 290
rect 290 288 292 290
rect 295 288 297 290
rect 3 278 5 280
rect 8 278 10 280
rect 13 278 15 280
rect 18 278 20 280
rect 23 278 25 280
rect 28 278 30 280
rect 33 278 35 280
rect 38 278 40 280
rect 43 278 45 280
rect 48 278 50 280
rect 53 278 55 280
rect 58 278 60 280
rect 63 278 65 280
rect 68 278 70 280
rect 73 278 75 280
rect 78 278 80 280
rect 83 278 85 280
rect 88 278 90 280
rect 93 278 95 280
rect 144 278 146 280
rect 149 278 151 280
rect 154 278 156 280
rect 205 278 207 280
rect 210 278 212 280
rect 215 278 217 280
rect 220 278 222 280
rect 225 278 227 280
rect 230 278 232 280
rect 235 278 237 280
rect 240 278 242 280
rect 245 278 247 280
rect 250 278 252 280
rect 255 278 257 280
rect 260 278 262 280
rect 265 278 267 280
rect 270 278 272 280
rect 275 278 277 280
rect 280 278 282 280
rect 285 278 287 280
rect 290 278 292 280
rect 295 278 297 280
rect 3 268 5 270
rect 8 268 10 270
rect 13 268 15 270
rect 18 268 20 270
rect 23 268 25 270
rect 28 268 30 270
rect 33 268 35 270
rect 38 268 40 270
rect 43 268 45 270
rect 48 268 50 270
rect 53 268 55 270
rect 58 268 60 270
rect 63 268 65 270
rect 68 268 70 270
rect 73 268 75 270
rect 78 268 80 270
rect 83 268 85 270
rect 88 268 90 270
rect 93 268 95 270
rect 144 268 146 270
rect 149 268 151 270
rect 154 268 156 270
rect 205 268 207 270
rect 210 268 212 270
rect 215 268 217 270
rect 220 268 222 270
rect 225 268 227 270
rect 230 268 232 270
rect 235 268 237 270
rect 240 268 242 270
rect 245 268 247 270
rect 250 268 252 270
rect 255 268 257 270
rect 260 268 262 270
rect 265 268 267 270
rect 270 268 272 270
rect 275 268 277 270
rect 280 268 282 270
rect 285 268 287 270
rect 290 268 292 270
rect 295 268 297 270
rect 8 258 10 260
rect 13 258 15 260
rect 18 258 20 260
rect 23 258 25 260
rect 28 258 30 260
rect 33 258 35 260
rect 38 258 40 260
rect 43 258 45 260
rect 48 258 50 260
rect 53 258 55 260
rect 58 258 60 260
rect 63 258 65 260
rect 68 258 70 260
rect 73 258 75 260
rect 78 258 80 260
rect 83 258 85 260
rect 88 258 90 260
rect 93 258 95 260
rect 144 258 146 260
rect 149 258 151 260
rect 154 258 156 260
rect 204 258 206 260
rect 209 258 211 260
rect 214 258 216 260
rect 219 258 221 260
rect 224 258 226 260
rect 229 258 231 260
rect 234 258 236 260
rect 239 258 241 260
rect 244 258 246 260
rect 249 258 251 260
rect 254 258 256 260
rect 259 258 261 260
rect 264 258 266 260
rect 269 258 271 260
rect 274 258 276 260
rect 279 258 281 260
rect 284 258 286 260
rect 289 258 291 260
rect 16 221 18 223
rect 21 221 23 223
rect 26 221 28 223
rect 31 221 33 223
rect 36 221 38 223
rect 41 221 43 223
rect 46 221 48 223
rect 51 221 53 223
rect 56 221 58 223
rect 61 221 63 223
rect 66 221 68 223
rect 71 221 73 223
rect 76 221 78 223
rect 81 221 83 223
rect 86 221 88 223
rect 91 221 93 223
rect 96 221 98 223
rect 101 221 103 223
rect 106 221 108 223
rect 111 221 113 223
rect 116 221 118 223
rect 121 221 123 223
rect 126 221 128 223
rect 131 221 133 223
rect 136 221 138 223
rect 141 221 143 223
rect 146 221 148 223
rect 151 221 153 223
rect 156 221 158 223
rect 161 221 163 223
rect 166 221 168 223
rect 171 221 173 223
rect 176 221 178 223
rect 181 221 183 223
rect 186 221 188 223
rect 191 221 193 223
rect 196 221 198 223
rect 201 221 203 223
rect 206 221 208 223
rect 211 221 213 223
rect 216 221 218 223
rect 221 221 223 223
rect 226 221 228 223
rect 231 221 233 223
rect 236 221 238 223
rect 241 221 243 223
rect 246 221 248 223
rect 251 221 253 223
rect 256 221 258 223
rect 261 221 263 223
rect 266 221 268 223
rect 271 221 273 223
rect 276 221 278 223
rect 281 221 283 223
rect 16 211 18 213
rect 21 211 23 213
rect 26 211 28 213
rect 31 211 33 213
rect 36 211 38 213
rect 41 211 43 213
rect 46 211 48 213
rect 51 211 53 213
rect 56 211 58 213
rect 61 211 63 213
rect 66 211 68 213
rect 71 211 73 213
rect 76 211 78 213
rect 81 211 83 213
rect 86 211 88 213
rect 91 211 93 213
rect 96 211 98 213
rect 101 211 103 213
rect 106 211 108 213
rect 111 211 113 213
rect 116 211 118 213
rect 121 211 123 213
rect 126 211 128 213
rect 131 211 133 213
rect 136 211 138 213
rect 141 211 143 213
rect 146 211 148 213
rect 151 211 153 213
rect 156 211 158 213
rect 161 211 163 213
rect 166 211 168 213
rect 171 211 173 213
rect 176 211 178 213
rect 181 211 183 213
rect 186 211 188 213
rect 191 211 193 213
rect 196 211 198 213
rect 201 211 203 213
rect 206 211 208 213
rect 211 211 213 213
rect 216 211 218 213
rect 221 211 223 213
rect 226 211 228 213
rect 231 211 233 213
rect 236 211 238 213
rect 241 211 243 213
rect 246 211 248 213
rect 251 211 253 213
rect 256 211 258 213
rect 261 211 263 213
rect 266 211 268 213
rect 271 211 273 213
rect 276 211 278 213
rect 281 211 283 213
rect 16 201 18 203
rect 21 201 23 203
rect 26 201 28 203
rect 31 201 33 203
rect 36 201 38 203
rect 41 201 43 203
rect 46 201 48 203
rect 51 201 53 203
rect 56 201 58 203
rect 61 201 63 203
rect 66 201 68 203
rect 71 201 73 203
rect 76 201 78 203
rect 81 201 83 203
rect 86 201 88 203
rect 91 201 93 203
rect 96 201 98 203
rect 101 201 103 203
rect 106 201 108 203
rect 111 201 113 203
rect 116 201 118 203
rect 121 201 123 203
rect 126 201 128 203
rect 131 201 133 203
rect 136 201 138 203
rect 141 201 143 203
rect 146 201 148 203
rect 151 201 153 203
rect 156 201 158 203
rect 161 201 163 203
rect 166 201 168 203
rect 171 201 173 203
rect 176 201 178 203
rect 181 201 183 203
rect 186 201 188 203
rect 191 201 193 203
rect 196 201 198 203
rect 201 201 203 203
rect 206 201 208 203
rect 211 201 213 203
rect 216 201 218 203
rect 221 201 223 203
rect 226 201 228 203
rect 231 201 233 203
rect 236 201 238 203
rect 241 201 243 203
rect 246 201 248 203
rect 251 201 253 203
rect 256 201 258 203
rect 261 201 263 203
rect 266 201 268 203
rect 271 201 273 203
rect 276 201 278 203
rect 281 201 283 203
rect 16 191 18 193
rect 21 191 23 193
rect 26 191 28 193
rect 31 191 33 193
rect 36 191 38 193
rect 41 191 43 193
rect 46 191 48 193
rect 51 191 53 193
rect 56 191 58 193
rect 61 191 63 193
rect 66 191 68 193
rect 71 191 73 193
rect 76 191 78 193
rect 81 191 83 193
rect 86 191 88 193
rect 91 191 93 193
rect 96 191 98 193
rect 101 191 103 193
rect 106 191 108 193
rect 111 191 113 193
rect 116 191 118 193
rect 121 191 123 193
rect 126 191 128 193
rect 131 191 133 193
rect 136 191 138 193
rect 141 191 143 193
rect 146 191 148 193
rect 151 191 153 193
rect 156 191 158 193
rect 161 191 163 193
rect 166 191 168 193
rect 171 191 173 193
rect 176 191 178 193
rect 181 191 183 193
rect 186 191 188 193
rect 191 191 193 193
rect 196 191 198 193
rect 201 191 203 193
rect 206 191 208 193
rect 211 191 213 193
rect 216 191 218 193
rect 221 191 223 193
rect 226 191 228 193
rect 231 191 233 193
rect 236 191 238 193
rect 241 191 243 193
rect 246 191 248 193
rect 251 191 253 193
rect 256 191 258 193
rect 261 191 263 193
rect 266 191 268 193
rect 271 191 273 193
rect 276 191 278 193
rect 281 191 283 193
rect 16 181 18 183
rect 21 181 23 183
rect 26 181 28 183
rect 31 181 33 183
rect 36 181 38 183
rect 41 181 43 183
rect 46 181 48 183
rect 51 181 53 183
rect 56 181 58 183
rect 61 181 63 183
rect 66 181 68 183
rect 71 181 73 183
rect 76 181 78 183
rect 81 181 83 183
rect 86 181 88 183
rect 91 181 93 183
rect 96 181 98 183
rect 101 181 103 183
rect 106 181 108 183
rect 111 181 113 183
rect 116 181 118 183
rect 121 181 123 183
rect 126 181 128 183
rect 131 181 133 183
rect 136 181 138 183
rect 141 181 143 183
rect 146 181 148 183
rect 151 181 153 183
rect 156 181 158 183
rect 161 181 163 183
rect 166 181 168 183
rect 171 181 173 183
rect 176 181 178 183
rect 181 181 183 183
rect 186 181 188 183
rect 191 181 193 183
rect 196 181 198 183
rect 201 181 203 183
rect 206 181 208 183
rect 211 181 213 183
rect 216 181 218 183
rect 221 181 223 183
rect 226 181 228 183
rect 231 181 233 183
rect 236 181 238 183
rect 241 181 243 183
rect 246 181 248 183
rect 251 181 253 183
rect 256 181 258 183
rect 261 181 263 183
rect 266 181 268 183
rect 271 181 273 183
rect 276 181 278 183
rect 281 181 283 183
rect 16 171 18 173
rect 21 171 23 173
rect 26 171 28 173
rect 31 171 33 173
rect 36 171 38 173
rect 41 171 43 173
rect 46 171 48 173
rect 51 171 53 173
rect 56 171 58 173
rect 61 171 63 173
rect 66 171 68 173
rect 71 171 73 173
rect 76 171 78 173
rect 81 171 83 173
rect 86 171 88 173
rect 91 171 93 173
rect 96 171 98 173
rect 101 171 103 173
rect 106 171 108 173
rect 111 171 113 173
rect 116 171 118 173
rect 121 171 123 173
rect 126 171 128 173
rect 131 171 133 173
rect 136 171 138 173
rect 141 171 143 173
rect 146 171 148 173
rect 151 171 153 173
rect 156 171 158 173
rect 161 171 163 173
rect 166 171 168 173
rect 171 171 173 173
rect 176 171 178 173
rect 181 171 183 173
rect 186 171 188 173
rect 191 171 193 173
rect 196 171 198 173
rect 201 171 203 173
rect 206 171 208 173
rect 211 171 213 173
rect 216 171 218 173
rect 221 171 223 173
rect 226 171 228 173
rect 231 171 233 173
rect 236 171 238 173
rect 241 171 243 173
rect 246 171 248 173
rect 251 171 253 173
rect 256 171 258 173
rect 261 171 263 173
rect 266 171 268 173
rect 271 171 273 173
rect 276 171 278 173
rect 281 171 283 173
rect 16 161 18 163
rect 21 161 23 163
rect 26 161 28 163
rect 31 161 33 163
rect 36 161 38 163
rect 41 161 43 163
rect 46 161 48 163
rect 51 161 53 163
rect 56 161 58 163
rect 61 161 63 163
rect 66 161 68 163
rect 71 161 73 163
rect 76 161 78 163
rect 81 161 83 163
rect 86 161 88 163
rect 91 161 93 163
rect 96 161 98 163
rect 101 161 103 163
rect 106 161 108 163
rect 111 161 113 163
rect 116 161 118 163
rect 121 161 123 163
rect 126 161 128 163
rect 131 161 133 163
rect 136 161 138 163
rect 141 161 143 163
rect 146 161 148 163
rect 151 161 153 163
rect 156 161 158 163
rect 161 161 163 163
rect 166 161 168 163
rect 171 161 173 163
rect 176 161 178 163
rect 181 161 183 163
rect 186 161 188 163
rect 191 161 193 163
rect 196 161 198 163
rect 201 161 203 163
rect 206 161 208 163
rect 211 161 213 163
rect 216 161 218 163
rect 221 161 223 163
rect 226 161 228 163
rect 231 161 233 163
rect 236 161 238 163
rect 241 161 243 163
rect 246 161 248 163
rect 251 161 253 163
rect 256 161 258 163
rect 261 161 263 163
rect 266 161 268 163
rect 271 161 273 163
rect 276 161 278 163
rect 281 161 283 163
rect 16 151 18 153
rect 21 151 23 153
rect 26 151 28 153
rect 31 151 33 153
rect 36 151 38 153
rect 41 151 43 153
rect 46 151 48 153
rect 51 151 53 153
rect 56 151 58 153
rect 61 151 63 153
rect 66 151 68 153
rect 71 151 73 153
rect 76 151 78 153
rect 81 151 83 153
rect 86 151 88 153
rect 91 151 93 153
rect 96 151 98 153
rect 101 151 103 153
rect 106 151 108 153
rect 111 151 113 153
rect 116 151 118 153
rect 121 151 123 153
rect 126 151 128 153
rect 131 151 133 153
rect 136 151 138 153
rect 141 151 143 153
rect 146 151 148 153
rect 151 151 153 153
rect 156 151 158 153
rect 161 151 163 153
rect 166 151 168 153
rect 171 151 173 153
rect 176 151 178 153
rect 181 151 183 153
rect 186 151 188 153
rect 191 151 193 153
rect 196 151 198 153
rect 201 151 203 153
rect 206 151 208 153
rect 211 151 213 153
rect 216 151 218 153
rect 221 151 223 153
rect 226 151 228 153
rect 231 151 233 153
rect 236 151 238 153
rect 241 151 243 153
rect 246 151 248 153
rect 251 151 253 153
rect 256 151 258 153
rect 261 151 263 153
rect 266 151 268 153
rect 271 151 273 153
rect 276 151 278 153
rect 281 151 283 153
rect 16 141 18 143
rect 21 141 23 143
rect 26 141 28 143
rect 31 141 33 143
rect 36 141 38 143
rect 41 141 43 143
rect 46 141 48 143
rect 51 141 53 143
rect 56 141 58 143
rect 61 141 63 143
rect 66 141 68 143
rect 71 141 73 143
rect 76 141 78 143
rect 81 141 83 143
rect 86 141 88 143
rect 91 141 93 143
rect 96 141 98 143
rect 101 141 103 143
rect 106 141 108 143
rect 111 141 113 143
rect 116 141 118 143
rect 121 141 123 143
rect 126 141 128 143
rect 131 141 133 143
rect 136 141 138 143
rect 141 141 143 143
rect 146 141 148 143
rect 151 141 153 143
rect 156 141 158 143
rect 161 141 163 143
rect 166 141 168 143
rect 171 141 173 143
rect 176 141 178 143
rect 181 141 183 143
rect 186 141 188 143
rect 191 141 193 143
rect 196 141 198 143
rect 201 141 203 143
rect 206 141 208 143
rect 211 141 213 143
rect 216 141 218 143
rect 221 141 223 143
rect 226 141 228 143
rect 231 141 233 143
rect 236 141 238 143
rect 241 141 243 143
rect 246 141 248 143
rect 251 141 253 143
rect 256 141 258 143
rect 261 141 263 143
rect 266 141 268 143
rect 271 141 273 143
rect 276 141 278 143
rect 281 141 283 143
rect 16 131 18 133
rect 21 131 23 133
rect 26 131 28 133
rect 31 131 33 133
rect 36 131 38 133
rect 41 131 43 133
rect 46 131 48 133
rect 51 131 53 133
rect 56 131 58 133
rect 61 131 63 133
rect 66 131 68 133
rect 71 131 73 133
rect 76 131 78 133
rect 81 131 83 133
rect 86 131 88 133
rect 91 131 93 133
rect 96 131 98 133
rect 101 131 103 133
rect 106 131 108 133
rect 111 131 113 133
rect 116 131 118 133
rect 121 131 123 133
rect 126 131 128 133
rect 131 131 133 133
rect 136 131 138 133
rect 141 131 143 133
rect 146 131 148 133
rect 151 131 153 133
rect 156 131 158 133
rect 161 131 163 133
rect 166 131 168 133
rect 171 131 173 133
rect 176 131 178 133
rect 181 131 183 133
rect 186 131 188 133
rect 191 131 193 133
rect 196 131 198 133
rect 201 131 203 133
rect 206 131 208 133
rect 211 131 213 133
rect 216 131 218 133
rect 221 131 223 133
rect 226 131 228 133
rect 231 131 233 133
rect 236 131 238 133
rect 241 131 243 133
rect 246 131 248 133
rect 251 131 253 133
rect 256 131 258 133
rect 261 131 263 133
rect 266 131 268 133
rect 271 131 273 133
rect 276 131 278 133
rect 281 131 283 133
rect 16 121 18 123
rect 21 121 23 123
rect 26 121 28 123
rect 31 121 33 123
rect 36 121 38 123
rect 41 121 43 123
rect 46 121 48 123
rect 51 121 53 123
rect 56 121 58 123
rect 61 121 63 123
rect 66 121 68 123
rect 71 121 73 123
rect 76 121 78 123
rect 81 121 83 123
rect 86 121 88 123
rect 91 121 93 123
rect 96 121 98 123
rect 101 121 103 123
rect 106 121 108 123
rect 111 121 113 123
rect 116 121 118 123
rect 121 121 123 123
rect 126 121 128 123
rect 131 121 133 123
rect 136 121 138 123
rect 141 121 143 123
rect 146 121 148 123
rect 151 121 153 123
rect 156 121 158 123
rect 161 121 163 123
rect 166 121 168 123
rect 171 121 173 123
rect 176 121 178 123
rect 181 121 183 123
rect 186 121 188 123
rect 191 121 193 123
rect 196 121 198 123
rect 201 121 203 123
rect 206 121 208 123
rect 211 121 213 123
rect 216 121 218 123
rect 221 121 223 123
rect 226 121 228 123
rect 231 121 233 123
rect 236 121 238 123
rect 241 121 243 123
rect 246 121 248 123
rect 251 121 253 123
rect 256 121 258 123
rect 261 121 263 123
rect 266 121 268 123
rect 271 121 273 123
rect 276 121 278 123
rect 281 121 283 123
rect 16 111 18 113
rect 21 111 23 113
rect 26 111 28 113
rect 31 111 33 113
rect 36 111 38 113
rect 41 111 43 113
rect 46 111 48 113
rect 51 111 53 113
rect 56 111 58 113
rect 61 111 63 113
rect 66 111 68 113
rect 71 111 73 113
rect 76 111 78 113
rect 81 111 83 113
rect 86 111 88 113
rect 91 111 93 113
rect 96 111 98 113
rect 101 111 103 113
rect 106 111 108 113
rect 111 111 113 113
rect 116 111 118 113
rect 121 111 123 113
rect 126 111 128 113
rect 131 111 133 113
rect 136 111 138 113
rect 141 111 143 113
rect 146 111 148 113
rect 151 111 153 113
rect 156 111 158 113
rect 161 111 163 113
rect 166 111 168 113
rect 171 111 173 113
rect 176 111 178 113
rect 181 111 183 113
rect 186 111 188 113
rect 191 111 193 113
rect 196 111 198 113
rect 201 111 203 113
rect 206 111 208 113
rect 211 111 213 113
rect 216 111 218 113
rect 221 111 223 113
rect 226 111 228 113
rect 231 111 233 113
rect 236 111 238 113
rect 241 111 243 113
rect 246 111 248 113
rect 251 111 253 113
rect 256 111 258 113
rect 261 111 263 113
rect 266 111 268 113
rect 271 111 273 113
rect 276 111 278 113
rect 281 111 283 113
rect 16 101 18 103
rect 21 101 23 103
rect 26 101 28 103
rect 31 101 33 103
rect 36 101 38 103
rect 41 101 43 103
rect 46 101 48 103
rect 51 101 53 103
rect 56 101 58 103
rect 61 101 63 103
rect 66 101 68 103
rect 71 101 73 103
rect 76 101 78 103
rect 81 101 83 103
rect 86 101 88 103
rect 91 101 93 103
rect 96 101 98 103
rect 101 101 103 103
rect 106 101 108 103
rect 111 101 113 103
rect 116 101 118 103
rect 121 101 123 103
rect 126 101 128 103
rect 131 101 133 103
rect 136 101 138 103
rect 141 101 143 103
rect 146 101 148 103
rect 151 101 153 103
rect 156 101 158 103
rect 161 101 163 103
rect 166 101 168 103
rect 171 101 173 103
rect 176 101 178 103
rect 181 101 183 103
rect 186 101 188 103
rect 191 101 193 103
rect 196 101 198 103
rect 201 101 203 103
rect 206 101 208 103
rect 211 101 213 103
rect 216 101 218 103
rect 221 101 223 103
rect 226 101 228 103
rect 231 101 233 103
rect 236 101 238 103
rect 241 101 243 103
rect 246 101 248 103
rect 251 101 253 103
rect 256 101 258 103
rect 261 101 263 103
rect 266 101 268 103
rect 271 101 273 103
rect 276 101 278 103
rect 281 101 283 103
rect 16 91 18 93
rect 21 91 23 93
rect 26 91 28 93
rect 31 91 33 93
rect 36 91 38 93
rect 41 91 43 93
rect 46 91 48 93
rect 51 91 53 93
rect 56 91 58 93
rect 61 91 63 93
rect 66 91 68 93
rect 71 91 73 93
rect 76 91 78 93
rect 81 91 83 93
rect 86 91 88 93
rect 91 91 93 93
rect 96 91 98 93
rect 101 91 103 93
rect 106 91 108 93
rect 111 91 113 93
rect 116 91 118 93
rect 121 91 123 93
rect 126 91 128 93
rect 131 91 133 93
rect 136 91 138 93
rect 141 91 143 93
rect 146 91 148 93
rect 151 91 153 93
rect 156 91 158 93
rect 161 91 163 93
rect 166 91 168 93
rect 171 91 173 93
rect 176 91 178 93
rect 181 91 183 93
rect 186 91 188 93
rect 191 91 193 93
rect 196 91 198 93
rect 201 91 203 93
rect 206 91 208 93
rect 211 91 213 93
rect 216 91 218 93
rect 221 91 223 93
rect 226 91 228 93
rect 231 91 233 93
rect 236 91 238 93
rect 241 91 243 93
rect 246 91 248 93
rect 251 91 253 93
rect 256 91 258 93
rect 261 91 263 93
rect 266 91 268 93
rect 271 91 273 93
rect 276 91 278 93
rect 281 91 283 93
rect 16 81 18 83
rect 21 81 23 83
rect 26 81 28 83
rect 31 81 33 83
rect 36 81 38 83
rect 41 81 43 83
rect 46 81 48 83
rect 51 81 53 83
rect 56 81 58 83
rect 61 81 63 83
rect 66 81 68 83
rect 71 81 73 83
rect 76 81 78 83
rect 81 81 83 83
rect 86 81 88 83
rect 91 81 93 83
rect 96 81 98 83
rect 101 81 103 83
rect 106 81 108 83
rect 111 81 113 83
rect 116 81 118 83
rect 121 81 123 83
rect 126 81 128 83
rect 131 81 133 83
rect 136 81 138 83
rect 141 81 143 83
rect 146 81 148 83
rect 151 81 153 83
rect 156 81 158 83
rect 161 81 163 83
rect 166 81 168 83
rect 171 81 173 83
rect 176 81 178 83
rect 181 81 183 83
rect 186 81 188 83
rect 191 81 193 83
rect 196 81 198 83
rect 201 81 203 83
rect 206 81 208 83
rect 211 81 213 83
rect 216 81 218 83
rect 221 81 223 83
rect 226 81 228 83
rect 231 81 233 83
rect 236 81 238 83
rect 241 81 243 83
rect 246 81 248 83
rect 251 81 253 83
rect 256 81 258 83
rect 261 81 263 83
rect 266 81 268 83
rect 271 81 273 83
rect 276 81 278 83
rect 281 81 283 83
rect 16 71 18 73
rect 21 71 23 73
rect 26 71 28 73
rect 31 71 33 73
rect 36 71 38 73
rect 41 71 43 73
rect 46 71 48 73
rect 51 71 53 73
rect 56 71 58 73
rect 61 71 63 73
rect 66 71 68 73
rect 71 71 73 73
rect 76 71 78 73
rect 81 71 83 73
rect 86 71 88 73
rect 91 71 93 73
rect 96 71 98 73
rect 101 71 103 73
rect 106 71 108 73
rect 111 71 113 73
rect 116 71 118 73
rect 121 71 123 73
rect 126 71 128 73
rect 131 71 133 73
rect 136 71 138 73
rect 141 71 143 73
rect 146 71 148 73
rect 151 71 153 73
rect 156 71 158 73
rect 161 71 163 73
rect 166 71 168 73
rect 171 71 173 73
rect 176 71 178 73
rect 181 71 183 73
rect 186 71 188 73
rect 191 71 193 73
rect 196 71 198 73
rect 201 71 203 73
rect 206 71 208 73
rect 211 71 213 73
rect 216 71 218 73
rect 221 71 223 73
rect 226 71 228 73
rect 231 71 233 73
rect 236 71 238 73
rect 241 71 243 73
rect 246 71 248 73
rect 251 71 253 73
rect 256 71 258 73
rect 261 71 263 73
rect 266 71 268 73
rect 271 71 273 73
rect 276 71 278 73
rect 281 71 283 73
rect 16 61 18 63
rect 21 61 23 63
rect 26 61 28 63
rect 31 61 33 63
rect 36 61 38 63
rect 41 61 43 63
rect 46 61 48 63
rect 51 61 53 63
rect 56 61 58 63
rect 61 61 63 63
rect 66 61 68 63
rect 71 61 73 63
rect 76 61 78 63
rect 81 61 83 63
rect 86 61 88 63
rect 91 61 93 63
rect 96 61 98 63
rect 101 61 103 63
rect 106 61 108 63
rect 111 61 113 63
rect 116 61 118 63
rect 121 61 123 63
rect 126 61 128 63
rect 131 61 133 63
rect 136 61 138 63
rect 141 61 143 63
rect 146 61 148 63
rect 151 61 153 63
rect 156 61 158 63
rect 161 61 163 63
rect 166 61 168 63
rect 171 61 173 63
rect 176 61 178 63
rect 181 61 183 63
rect 186 61 188 63
rect 191 61 193 63
rect 196 61 198 63
rect 201 61 203 63
rect 206 61 208 63
rect 211 61 213 63
rect 216 61 218 63
rect 221 61 223 63
rect 226 61 228 63
rect 231 61 233 63
rect 236 61 238 63
rect 241 61 243 63
rect 246 61 248 63
rect 251 61 253 63
rect 256 61 258 63
rect 261 61 263 63
rect 266 61 268 63
rect 271 61 273 63
rect 276 61 278 63
rect 281 61 283 63
rect 16 51 18 53
rect 21 51 23 53
rect 26 51 28 53
rect 31 51 33 53
rect 36 51 38 53
rect 41 51 43 53
rect 46 51 48 53
rect 51 51 53 53
rect 56 51 58 53
rect 61 51 63 53
rect 66 51 68 53
rect 71 51 73 53
rect 76 51 78 53
rect 81 51 83 53
rect 86 51 88 53
rect 91 51 93 53
rect 96 51 98 53
rect 101 51 103 53
rect 106 51 108 53
rect 111 51 113 53
rect 116 51 118 53
rect 121 51 123 53
rect 126 51 128 53
rect 131 51 133 53
rect 136 51 138 53
rect 141 51 143 53
rect 146 51 148 53
rect 151 51 153 53
rect 156 51 158 53
rect 161 51 163 53
rect 166 51 168 53
rect 171 51 173 53
rect 176 51 178 53
rect 181 51 183 53
rect 186 51 188 53
rect 191 51 193 53
rect 196 51 198 53
rect 201 51 203 53
rect 206 51 208 53
rect 211 51 213 53
rect 216 51 218 53
rect 221 51 223 53
rect 226 51 228 53
rect 231 51 233 53
rect 236 51 238 53
rect 241 51 243 53
rect 246 51 248 53
rect 251 51 253 53
rect 256 51 258 53
rect 261 51 263 53
rect 266 51 268 53
rect 271 51 273 53
rect 276 51 278 53
rect 281 51 283 53
rect 16 41 18 43
rect 21 41 23 43
rect 26 41 28 43
rect 31 41 33 43
rect 36 41 38 43
rect 41 41 43 43
rect 46 41 48 43
rect 51 41 53 43
rect 56 41 58 43
rect 61 41 63 43
rect 66 41 68 43
rect 71 41 73 43
rect 76 41 78 43
rect 81 41 83 43
rect 86 41 88 43
rect 91 41 93 43
rect 96 41 98 43
rect 101 41 103 43
rect 106 41 108 43
rect 111 41 113 43
rect 116 41 118 43
rect 121 41 123 43
rect 126 41 128 43
rect 131 41 133 43
rect 136 41 138 43
rect 141 41 143 43
rect 146 41 148 43
rect 151 41 153 43
rect 156 41 158 43
rect 161 41 163 43
rect 166 41 168 43
rect 171 41 173 43
rect 176 41 178 43
rect 181 41 183 43
rect 186 41 188 43
rect 191 41 193 43
rect 196 41 198 43
rect 201 41 203 43
rect 206 41 208 43
rect 211 41 213 43
rect 216 41 218 43
rect 221 41 223 43
rect 226 41 228 43
rect 231 41 233 43
rect 236 41 238 43
rect 241 41 243 43
rect 246 41 248 43
rect 251 41 253 43
rect 256 41 258 43
rect 261 41 263 43
rect 266 41 268 43
rect 271 41 273 43
rect 276 41 278 43
rect 281 41 283 43
rect 16 31 18 33
rect 21 31 23 33
rect 26 31 28 33
rect 31 31 33 33
rect 36 31 38 33
rect 41 31 43 33
rect 46 31 48 33
rect 51 31 53 33
rect 56 31 58 33
rect 61 31 63 33
rect 66 31 68 33
rect 71 31 73 33
rect 76 31 78 33
rect 81 31 83 33
rect 86 31 88 33
rect 91 31 93 33
rect 96 31 98 33
rect 101 31 103 33
rect 106 31 108 33
rect 111 31 113 33
rect 116 31 118 33
rect 121 31 123 33
rect 126 31 128 33
rect 131 31 133 33
rect 136 31 138 33
rect 141 31 143 33
rect 146 31 148 33
rect 151 31 153 33
rect 156 31 158 33
rect 161 31 163 33
rect 166 31 168 33
rect 171 31 173 33
rect 176 31 178 33
rect 181 31 183 33
rect 186 31 188 33
rect 191 31 193 33
rect 196 31 198 33
rect 201 31 203 33
rect 206 31 208 33
rect 211 31 213 33
rect 216 31 218 33
rect 221 31 223 33
rect 226 31 228 33
rect 231 31 233 33
rect 236 31 238 33
rect 241 31 243 33
rect 246 31 248 33
rect 251 31 253 33
rect 256 31 258 33
rect 261 31 263 33
rect 266 31 268 33
rect 271 31 273 33
rect 276 31 278 33
rect 281 31 283 33
rect 16 21 18 23
rect 21 21 23 23
rect 26 21 28 23
rect 31 21 33 23
rect 36 21 38 23
rect 41 21 43 23
rect 46 21 48 23
rect 51 21 53 23
rect 56 21 58 23
rect 61 21 63 23
rect 66 21 68 23
rect 71 21 73 23
rect 76 21 78 23
rect 81 21 83 23
rect 86 21 88 23
rect 91 21 93 23
rect 96 21 98 23
rect 101 21 103 23
rect 106 21 108 23
rect 111 21 113 23
rect 116 21 118 23
rect 121 21 123 23
rect 126 21 128 23
rect 131 21 133 23
rect 136 21 138 23
rect 141 21 143 23
rect 146 21 148 23
rect 151 21 153 23
rect 156 21 158 23
rect 161 21 163 23
rect 166 21 168 23
rect 171 21 173 23
rect 176 21 178 23
rect 181 21 183 23
rect 186 21 188 23
rect 191 21 193 23
rect 196 21 198 23
rect 201 21 203 23
rect 206 21 208 23
rect 211 21 213 23
rect 216 21 218 23
rect 221 21 223 23
rect 226 21 228 23
rect 231 21 233 23
rect 236 21 238 23
rect 241 21 243 23
rect 246 21 248 23
rect 251 21 253 23
rect 256 21 258 23
rect 261 21 263 23
rect 266 21 268 23
rect 271 21 273 23
rect 276 21 278 23
rect 281 21 283 23
rect 104 3 106 5
rect 109 3 111 5
rect 114 3 116 5
rect 119 3 121 5
rect 124 3 126 5
rect 129 3 131 5
rect 134 3 136 5
rect 139 3 141 5
rect 144 3 146 5
rect 149 3 151 5
rect 154 3 156 5
rect 159 3 161 5
rect 164 3 166 5
rect 169 3 171 5
rect 174 3 176 5
rect 179 3 181 5
rect 184 3 186 5
rect 189 3 191 5
rect 194 3 196 5
<< metal3 >>
rect 23 743 277 997
<< gv2 >>
rect 47 971 49 973
rect 59 971 61 973
rect 71 971 73 973
rect 83 971 85 973
rect 95 971 97 973
rect 107 971 109 973
rect 119 971 121 973
rect 131 971 133 973
rect 143 971 145 973
rect 155 971 157 973
rect 167 971 169 973
rect 179 971 181 973
rect 191 971 193 973
rect 203 971 205 973
rect 215 971 217 973
rect 227 971 229 973
rect 239 971 241 973
rect 251 971 253 973
rect 47 959 49 961
rect 59 959 61 961
rect 71 959 73 961
rect 83 959 85 961
rect 95 959 97 961
rect 107 959 109 961
rect 119 959 121 961
rect 131 959 133 961
rect 143 959 145 961
rect 155 959 157 961
rect 167 959 169 961
rect 179 959 181 961
rect 191 959 193 961
rect 203 959 205 961
rect 215 959 217 961
rect 227 959 229 961
rect 239 959 241 961
rect 251 959 253 961
rect 47 947 49 949
rect 59 947 61 949
rect 71 947 73 949
rect 83 947 85 949
rect 95 947 97 949
rect 107 947 109 949
rect 119 947 121 949
rect 131 947 133 949
rect 143 947 145 949
rect 155 947 157 949
rect 167 947 169 949
rect 179 947 181 949
rect 191 947 193 949
rect 203 947 205 949
rect 215 947 217 949
rect 227 947 229 949
rect 239 947 241 949
rect 251 947 253 949
rect 47 935 49 937
rect 59 935 61 937
rect 71 935 73 937
rect 83 935 85 937
rect 95 935 97 937
rect 107 935 109 937
rect 119 935 121 937
rect 131 935 133 937
rect 143 935 145 937
rect 155 935 157 937
rect 167 935 169 937
rect 179 935 181 937
rect 191 935 193 937
rect 203 935 205 937
rect 215 935 217 937
rect 227 935 229 937
rect 239 935 241 937
rect 251 935 253 937
rect 47 923 49 925
rect 59 923 61 925
rect 71 923 73 925
rect 83 923 85 925
rect 95 923 97 925
rect 107 923 109 925
rect 119 923 121 925
rect 131 923 133 925
rect 143 923 145 925
rect 155 923 157 925
rect 167 923 169 925
rect 179 923 181 925
rect 191 923 193 925
rect 203 923 205 925
rect 215 923 217 925
rect 227 923 229 925
rect 239 923 241 925
rect 251 923 253 925
rect 47 911 49 913
rect 59 911 61 913
rect 71 911 73 913
rect 83 911 85 913
rect 95 911 97 913
rect 107 911 109 913
rect 119 911 121 913
rect 131 911 133 913
rect 143 911 145 913
rect 155 911 157 913
rect 167 911 169 913
rect 179 911 181 913
rect 191 911 193 913
rect 203 911 205 913
rect 215 911 217 913
rect 227 911 229 913
rect 239 911 241 913
rect 251 911 253 913
rect 47 899 49 901
rect 59 899 61 901
rect 71 899 73 901
rect 83 899 85 901
rect 95 899 97 901
rect 107 899 109 901
rect 119 899 121 901
rect 131 899 133 901
rect 143 899 145 901
rect 155 899 157 901
rect 167 899 169 901
rect 179 899 181 901
rect 191 899 193 901
rect 203 899 205 901
rect 215 899 217 901
rect 227 899 229 901
rect 239 899 241 901
rect 251 899 253 901
rect 47 887 49 889
rect 59 887 61 889
rect 71 887 73 889
rect 83 887 85 889
rect 95 887 97 889
rect 107 887 109 889
rect 119 887 121 889
rect 131 887 133 889
rect 143 887 145 889
rect 155 887 157 889
rect 167 887 169 889
rect 179 887 181 889
rect 191 887 193 889
rect 203 887 205 889
rect 215 887 217 889
rect 227 887 229 889
rect 239 887 241 889
rect 251 887 253 889
rect 47 875 49 877
rect 59 875 61 877
rect 71 875 73 877
rect 83 875 85 877
rect 95 875 97 877
rect 107 875 109 877
rect 119 875 121 877
rect 131 875 133 877
rect 143 875 145 877
rect 155 875 157 877
rect 167 875 169 877
rect 179 875 181 877
rect 191 875 193 877
rect 203 875 205 877
rect 215 875 217 877
rect 227 875 229 877
rect 239 875 241 877
rect 251 875 253 877
rect 47 863 49 865
rect 59 863 61 865
rect 71 863 73 865
rect 83 863 85 865
rect 95 863 97 865
rect 107 863 109 865
rect 119 863 121 865
rect 131 863 133 865
rect 143 863 145 865
rect 155 863 157 865
rect 167 863 169 865
rect 179 863 181 865
rect 191 863 193 865
rect 203 863 205 865
rect 215 863 217 865
rect 227 863 229 865
rect 239 863 241 865
rect 251 863 253 865
rect 47 851 49 853
rect 59 851 61 853
rect 71 851 73 853
rect 83 851 85 853
rect 95 851 97 853
rect 107 851 109 853
rect 119 851 121 853
rect 131 851 133 853
rect 143 851 145 853
rect 155 851 157 853
rect 167 851 169 853
rect 179 851 181 853
rect 191 851 193 853
rect 203 851 205 853
rect 215 851 217 853
rect 227 851 229 853
rect 239 851 241 853
rect 251 851 253 853
rect 47 839 49 841
rect 59 839 61 841
rect 71 839 73 841
rect 83 839 85 841
rect 95 839 97 841
rect 107 839 109 841
rect 119 839 121 841
rect 131 839 133 841
rect 143 839 145 841
rect 155 839 157 841
rect 167 839 169 841
rect 179 839 181 841
rect 191 839 193 841
rect 203 839 205 841
rect 215 839 217 841
rect 227 839 229 841
rect 239 839 241 841
rect 251 839 253 841
rect 47 827 49 829
rect 59 827 61 829
rect 71 827 73 829
rect 83 827 85 829
rect 95 827 97 829
rect 107 827 109 829
rect 119 827 121 829
rect 131 827 133 829
rect 143 827 145 829
rect 155 827 157 829
rect 167 827 169 829
rect 179 827 181 829
rect 191 827 193 829
rect 203 827 205 829
rect 215 827 217 829
rect 227 827 229 829
rect 239 827 241 829
rect 251 827 253 829
rect 47 815 49 817
rect 59 815 61 817
rect 71 815 73 817
rect 83 815 85 817
rect 95 815 97 817
rect 107 815 109 817
rect 119 815 121 817
rect 131 815 133 817
rect 143 815 145 817
rect 155 815 157 817
rect 167 815 169 817
rect 179 815 181 817
rect 191 815 193 817
rect 203 815 205 817
rect 215 815 217 817
rect 227 815 229 817
rect 239 815 241 817
rect 251 815 253 817
rect 47 803 49 805
rect 59 803 61 805
rect 71 803 73 805
rect 83 803 85 805
rect 95 803 97 805
rect 107 803 109 805
rect 119 803 121 805
rect 131 803 133 805
rect 143 803 145 805
rect 155 803 157 805
rect 167 803 169 805
rect 179 803 181 805
rect 191 803 193 805
rect 203 803 205 805
rect 215 803 217 805
rect 227 803 229 805
rect 239 803 241 805
rect 251 803 253 805
rect 47 791 49 793
rect 59 791 61 793
rect 71 791 73 793
rect 83 791 85 793
rect 95 791 97 793
rect 107 791 109 793
rect 119 791 121 793
rect 131 791 133 793
rect 143 791 145 793
rect 155 791 157 793
rect 167 791 169 793
rect 179 791 181 793
rect 191 791 193 793
rect 203 791 205 793
rect 215 791 217 793
rect 227 791 229 793
rect 239 791 241 793
rect 251 791 253 793
rect 47 779 49 781
rect 59 779 61 781
rect 71 779 73 781
rect 83 779 85 781
rect 95 779 97 781
rect 107 779 109 781
rect 119 779 121 781
rect 131 779 133 781
rect 143 779 145 781
rect 155 779 157 781
rect 167 779 169 781
rect 179 779 181 781
rect 191 779 193 781
rect 203 779 205 781
rect 215 779 217 781
rect 227 779 229 781
rect 239 779 241 781
rect 251 779 253 781
rect 47 767 49 769
rect 59 767 61 769
rect 71 767 73 769
rect 83 767 85 769
rect 95 767 97 769
rect 107 767 109 769
rect 119 767 121 769
rect 131 767 133 769
rect 143 767 145 769
rect 155 767 157 769
rect 167 767 169 769
rect 179 767 181 769
rect 191 767 193 769
rect 203 767 205 769
rect 215 767 217 769
rect 227 767 229 769
rect 239 767 241 769
rect 251 767 253 769
<< glass >>
rect 43 763 257 977
<< xp >>
rect 23 743 277 997
<< labels >>
rlabel metal1 150 0 150 0 8 GND!
rlabel metal2 132 540 132 540 6 vdd:2
rlabel metal1 150 -8 150 -8 8 GND!
<< end >>
