magic
tech scmos
timestamp 1683038052
<< metal1 >>
rect -2 -2 2 2
<< metal2 >>
rect -2 -2 2 2
<< gv1 >>
rect -1 -1 1 1
<< end >>
