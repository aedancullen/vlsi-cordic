magic
tech scmos
timestamp 1683038052
<< polysilicon >>
rect 2084 3345 3264 3346
rect 2084 3159 3269 3345
rect 2084 3043 3032 3159
rect 1051 3040 3032 3043
rect 1051 2799 3031 3040
rect 1021 1818 3192 2728
rect -909 -1143 -216 1021
rect -85 -755 870 1015
rect 985 -703 3249 1681
rect 2476 -1359 3249 -703
<< metal1 >>
rect -1375 4088 -1314 4128
rect -1080 4097 -1019 4137
rect -778 4096 -717 4136
rect -482 4096 -421 4136
rect -170 4093 -109 4133
rect 121 4085 182 4125
rect 421 4086 470 4129
rect 715 4093 776 4133
rect 1023 4093 1084 4133
rect 1311 4085 1372 4125
rect 1621 4093 1682 4133
rect 1915 4085 1976 4125
rect -2232 3222 -2190 3282
rect -2230 2916 -2188 2976
rect 399 2740 498 3389
rect 2084 3345 3264 3346
rect 918 3236 924 3304
rect 930 3236 936 3320
rect 942 3236 948 3288
rect 978 3107 984 3320
rect 990 3107 996 3263
rect 1315 3207 1408 3215
rect 2084 3159 3269 3345
rect 3981 3228 4021 3269
rect 2084 3043 3032 3159
rect 1051 3040 3032 3043
rect 894 2857 1020 2864
rect 1051 2799 3031 3040
rect 3992 2934 4032 2975
rect 3288 2910 3292 2915
rect -2230 2629 -2188 2689
rect -2232 2326 -2190 2386
rect -1491 2179 -945 2180
rect -1491 2099 -823 2179
rect -1491 2095 -945 2099
rect -2229 2021 -2189 2083
rect -1492 2060 -945 2095
rect -1492 2040 -1019 2060
rect -891 2051 -879 2056
rect 894 2051 900 2056
rect -1492 2004 -1455 2040
rect 894 2031 900 2037
rect -954 2011 -913 2016
rect 894 2011 900 2016
rect 894 1991 900 1996
rect 894 1971 900 1976
rect -892 1921 -879 1926
rect 1021 1818 3192 2728
rect 3994 2641 4034 2682
rect 3285 2611 3289 2616
rect 3288 2311 3292 2315
rect -892 1811 -879 1816
rect 894 1811 900 1816
rect -2233 1716 -2191 1776
rect 821 1709 3293 1796
rect 824 1708 3289 1709
rect -892 1691 -879 1696
rect -892 1491 -870 1496
rect -2232 1425 -2190 1485
rect -891 1291 -873 1296
rect -892 1241 -874 1246
rect -2229 1116 -2187 1176
rect -2229 825 -2187 885
rect -2226 523 -2184 583
rect -2235 -78 -2193 -18
rect -2228 -382 -2186 -322
rect -2229 -679 -2187 -619
rect -1493 -689 -1488 -685
rect -2225 -977 -2183 -917
rect -1491 -989 -1487 -985
rect -909 -1143 -216 1021
rect -1494 -1289 -1488 -1285
rect -1389 -1393 -1385 -1387
rect -1089 -1392 -1085 -1386
rect -789 -1394 -785 -1388
rect -198 -1392 -97 1048
rect -85 -755 870 1015
rect 985 -703 3249 1681
rect 2476 -1359 3249 -703
rect 111 -1374 115 -1372
rect 22 -1378 115 -1374
rect 22 -1386 26 -1378
rect 111 -1390 115 -1378
rect 411 -1391 415 -1385
rect 711 -1394 715 -1388
rect 1011 -1393 1015 -1387
rect 1311 -1394 1315 -1388
rect 1910 -1395 1914 -1389
rect 2210 -1393 2214 -1387
rect -1077 -2134 -1029 -2092
rect -774 -2129 -726 -2087
rect -476 -2127 -428 -2085
rect 118 -2130 166 -2088
rect 429 -2130 477 -2088
rect 732 -2130 780 -2088
rect 1033 -2125 1081 -2083
rect 1331 -2127 1379 -2085
rect 1927 -2133 1975 -2091
rect 2231 -2136 2279 -2094
rect 2523 -2130 2571 -2088
<< metal2 >>
rect -1477 3378 -1471 3381
rect -1405 3378 -1399 3392
rect -1241 3379 -1234 3384
rect -1477 3372 -1399 3378
rect -1177 3368 -1171 3381
rect -1103 3368 -1097 3392
rect -940 3381 -936 3385
rect -1488 3359 -1484 3363
rect -1177 3362 -1097 3368
rect -877 3366 -871 3381
rect -805 3366 -799 3391
rect -640 3381 -636 3385
rect -877 3360 -799 3366
rect -577 3368 -571 3381
rect -506 3368 -500 3392
rect -339 3381 -335 3385
rect -577 3362 -500 3368
rect -277 3368 -271 3381
rect -204 3368 -198 3391
rect -39 3381 -35 3385
rect 23 3374 29 3381
rect 95 3374 101 3392
rect 261 3382 265 3387
rect 23 3368 101 3374
rect 623 3369 629 3381
rect 694 3369 700 3392
rect 861 3381 865 3385
rect -277 3362 -198 3368
rect 623 3363 700 3369
rect 923 3370 929 3381
rect 995 3370 1001 3392
rect 1160 3381 1164 3385
rect 923 3364 1001 3370
rect 1223 3371 1229 3381
rect 1293 3371 1299 3391
rect 1459 3380 1463 3384
rect 1223 3365 1299 3371
rect 1523 3366 1529 3381
rect 1597 3366 1603 3392
rect 1760 3381 1764 3385
rect 1523 3360 1603 3366
rect 1823 3360 1829 3381
rect 1896 3360 1902 3392
rect 2057 3380 2061 3384
rect 2123 3376 2127 3386
rect 2195 3376 2199 3389
rect 2123 3372 2199 3376
rect 2723 3375 2727 3385
rect 2795 3375 2799 3388
rect 2723 3371 2799 3375
rect 3024 3377 3028 3383
rect 3095 3377 3099 3388
rect 3024 3373 3099 3377
rect 1823 3354 1902 3360
rect 2084 3345 3264 3346
rect 918 3236 924 3304
rect 930 3236 936 3320
rect 942 3236 948 3288
rect -1493 3193 -1467 3199
rect -1473 3129 -1467 3193
rect -1481 3123 -1467 3129
rect 978 3107 984 3320
rect 990 3107 996 3263
rect 1315 3207 1408 3215
rect 2084 3159 3269 3345
rect -1481 3057 -1433 3066
rect -1445 3056 -1434 3057
rect 2084 3043 3032 3159
rect 1051 3040 3032 3043
rect 3062 3149 3287 3152
rect -1492 2894 -1463 2900
rect -1469 2829 -1463 2894
rect 894 2857 1020 2864
rect -1482 2823 -1463 2829
rect 1051 2799 3031 3040
rect 3062 2791 3065 3149
rect 3259 3123 3281 3129
rect 3259 2915 3265 3123
rect 3259 2909 3292 2915
rect -442 2788 3065 2791
rect 3200 2849 3286 2852
rect -1481 2765 -1436 2766
rect -1481 2757 -1434 2765
rect -442 2761 -439 2788
rect 3200 2769 3203 2849
rect -150 2766 3203 2769
rect 3262 2823 3281 2829
rect -1445 2756 -1434 2757
rect -462 2752 -438 2761
rect -350 2752 -346 2756
rect -150 2755 -147 2766
rect 105 2756 3220 2761
rect -22 2752 -18 2756
rect 90 2752 94 2756
rect -1493 2594 -1467 2600
rect -1473 2529 -1467 2594
rect -1481 2523 -1467 2529
rect -1481 2457 -1434 2466
rect -1445 2456 -1434 2457
rect -1494 2296 -1462 2302
rect -1468 2229 -1462 2296
rect -1481 2223 -1462 2229
rect -839 2101 -824 2177
rect -1000 2052 -881 2056
rect 890 2052 972 2056
rect -1000 2051 -885 2052
rect 894 2051 972 2052
rect -1481 1871 -1468 1877
rect -1474 1807 -1468 1871
rect -1492 1801 -1468 1807
rect -1481 1642 -1435 1643
rect -1481 1634 -1434 1642
rect -1445 1633 -1434 1634
rect -1481 1565 -1435 1566
rect -1481 1557 -1434 1565
rect -1445 1556 -1434 1557
rect -1492 1393 -1465 1399
rect -1471 1329 -1465 1393
rect -1481 1323 -1465 1329
rect -1481 1257 -1434 1266
rect -1445 1256 -1434 1257
rect -1494 1093 -1464 1099
rect -1470 1029 -1464 1093
rect -1481 1023 -1464 1029
rect -1481 957 -1434 966
rect -1445 956 -1434 957
rect -1490 792 -1463 798
rect -1469 729 -1463 792
rect -1481 723 -1463 729
rect -1481 657 -1434 666
rect -1445 656 -1434 657
rect -1493 495 -1462 501
rect -1468 429 -1462 495
rect -1481 423 -1462 429
rect -1481 71 -1450 77
rect -1456 5 -1450 71
rect -1492 -1 -1450 5
rect -1489 -164 -1482 -159
rect -1000 -448 -994 2051
rect 894 2036 960 2037
rect 890 2032 960 2036
rect 894 2031 960 2032
rect -954 2012 -946 2016
rect -928 2012 -920 2016
rect 890 2012 948 2016
rect 894 2011 948 2012
rect 890 1992 936 1996
rect 894 1991 936 1992
rect 890 1972 924 1976
rect 894 1971 924 1972
rect -1490 -454 -994 -448
rect -988 1925 -892 1926
rect -988 1921 -884 1925
rect -1481 -477 -1463 -471
rect -1469 -684 -1463 -477
rect -1493 -690 -1463 -684
rect -988 -749 -982 1921
rect -1488 -755 -982 -749
rect -976 1815 -892 1816
rect -976 1811 -884 1815
rect 890 1812 912 1816
rect 894 1811 912 1812
rect -1481 -777 -1454 -771
rect -1460 -984 -1454 -777
rect -1492 -990 -1454 -984
rect -976 -1049 -970 1811
rect 890 1792 900 1796
rect 827 1709 844 1784
rect -1485 -1055 -970 -1049
rect -964 1695 -892 1696
rect -964 1691 -884 1695
rect -1481 -1077 -1465 -1071
rect -1471 -1284 -1465 -1077
rect -964 -1144 -958 1691
rect -1494 -1290 -1465 -1284
rect -1151 -1150 -958 -1144
rect -952 1495 -892 1496
rect -952 1491 -884 1495
rect -1492 -1308 -1471 -1302
rect -1477 -1371 -1471 -1308
rect -1390 -1371 -1171 -1365
rect -1485 -1377 -1470 -1371
rect -1477 -1381 -1471 -1377
rect -1390 -1393 -1384 -1371
rect -1177 -1381 -1171 -1371
rect -1151 -1389 -1145 -1150
rect -952 -1224 -946 1491
rect -940 1295 -891 1296
rect -940 1291 -883 1295
rect -940 -1191 -934 1291
rect -928 1245 -892 1246
rect -928 1241 -884 1245
rect -928 -1157 -922 1241
rect -909 -1143 -216 1021
rect -85 -755 870 1015
rect 894 -767 900 1792
rect 346 -773 900 -767
rect -928 -1163 47 -1157
rect -940 -1197 -555 -1191
rect -952 -1230 -844 -1224
rect -1091 -1374 -871 -1368
rect -1091 -1392 -1085 -1374
rect -877 -1382 -871 -1374
rect -850 -1384 -844 -1230
rect -791 -1377 -571 -1371
rect -791 -1394 -785 -1377
rect -577 -1381 -571 -1377
rect -561 -1382 -555 -1197
rect -561 -1388 -549 -1382
rect 22 -1386 26 -1380
rect 41 -1391 47 -1163
rect 323 -1370 329 -1369
rect 109 -1376 329 -1370
rect 110 -1378 116 -1376
rect 323 -1381 329 -1376
rect 346 -1390 352 -773
rect 906 -802 912 1811
rect 639 -808 912 -802
rect 410 -1374 629 -1368
rect 410 -1392 416 -1374
rect 623 -1381 629 -1374
rect 639 -1384 645 -808
rect 918 -848 924 1971
rect 930 -817 936 1991
rect 942 -787 948 2011
rect 954 -755 960 2031
rect 966 -716 972 2051
rect 1021 1818 3192 2728
rect 3215 2551 3220 2756
rect 3262 2616 3268 2823
rect 3262 2610 3289 2616
rect 3215 2546 3286 2551
rect 3257 2523 3281 2529
rect 3257 2317 3263 2523
rect 3257 2311 3292 2317
rect 3266 2295 3289 2299
rect 3266 2228 3270 2295
rect 3266 2224 3286 2228
rect 3266 1995 3288 1999
rect 3266 1930 3270 1995
rect 3266 1926 3286 1930
rect 985 -703 3249 1681
rect 3271 1395 3289 1399
rect 3271 1329 3275 1395
rect 3271 1325 3286 1329
rect 3273 1095 3288 1099
rect 3273 1028 3277 1095
rect 3273 1024 3288 1028
rect 3269 795 3289 799
rect 3269 729 3273 795
rect 3269 725 3286 729
rect 3269 495 3289 499
rect 3269 429 3273 495
rect 3269 425 3285 429
rect 3269 195 3290 199
rect 3269 128 3273 195
rect 3269 124 3286 128
rect 3270 -405 3288 -401
rect 3270 -473 3274 -405
rect 3270 -477 3285 -473
rect 966 -722 2450 -716
rect 954 -761 2148 -755
rect 942 -793 1848 -787
rect 930 -823 1263 -817
rect 918 -854 950 -848
rect 709 -1372 929 -1366
rect 709 -1394 715 -1372
rect 923 -1384 929 -1372
rect 944 -1386 950 -854
rect 1011 -1376 1229 -1370
rect 1011 -1393 1017 -1376
rect 1223 -1381 1229 -1376
rect 1243 -1392 1249 -823
rect 1310 -1368 1829 -1362
rect 1310 -1394 1316 -1368
rect 1823 -1381 1829 -1368
rect 1842 -1389 1848 -793
rect 1909 -1374 2129 -1368
rect 1909 -1397 1915 -1374
rect 2123 -1382 2129 -1374
rect 2142 -1387 2148 -761
rect 2208 -1365 2429 -1359
rect 2208 -1393 2214 -1365
rect 2423 -1382 2429 -1365
rect 2444 -1391 2450 -722
rect 2476 -1359 3249 -703
rect 3269 -705 3288 -701
rect 3269 -773 3273 -705
rect 3269 -777 3286 -773
rect 3270 -1005 3289 -1001
rect 3270 -1072 3274 -1005
rect 3270 -1076 3284 -1072
rect 3272 -1305 3288 -1301
rect 3272 -1372 3276 -1305
rect 2722 -1377 2799 -1373
rect 2722 -1384 2726 -1377
rect 2795 -1389 2799 -1377
rect 3024 -1377 3099 -1373
rect 3272 -1376 3286 -1372
rect 3024 -1388 3028 -1377
rect 3095 -1389 3099 -1377
<< gv1 >>
rect 3289 2911 3291 2913
rect 3286 2612 3288 2614
rect 3289 2312 3291 2314
rect -838 2173 -836 2175
rect -833 2173 -831 2175
rect -828 2173 -826 2175
rect -838 2168 -836 2170
rect -833 2168 -831 2170
rect -828 2168 -826 2170
rect -838 2163 -836 2165
rect -833 2163 -831 2165
rect -828 2163 -826 2165
rect -838 2158 -836 2160
rect -833 2158 -831 2160
rect -828 2158 -826 2160
rect -838 2153 -836 2155
rect -833 2153 -831 2155
rect -828 2153 -826 2155
rect -838 2148 -836 2150
rect -833 2148 -831 2150
rect -828 2148 -826 2150
rect -838 2143 -836 2145
rect -833 2143 -831 2145
rect -828 2143 -826 2145
rect -838 2138 -836 2140
rect -833 2138 -831 2140
rect -828 2138 -826 2140
rect -838 2133 -836 2135
rect -833 2133 -831 2135
rect -828 2133 -826 2135
rect -838 2128 -836 2130
rect -833 2128 -831 2130
rect -828 2128 -826 2130
rect -838 2123 -836 2125
rect -833 2123 -831 2125
rect -828 2123 -826 2125
rect -838 2118 -836 2120
rect -833 2118 -831 2120
rect -828 2118 -826 2120
rect -838 2113 -836 2115
rect -833 2113 -831 2115
rect -828 2113 -826 2115
rect -838 2108 -836 2110
rect -833 2108 -831 2110
rect -828 2108 -826 2110
rect -838 2103 -836 2105
rect -833 2103 -831 2105
rect -828 2103 -826 2105
rect -889 2052 -887 2054
rect 896 2052 898 2054
rect 896 2033 898 2035
rect -949 2013 -947 2015
rect -927 2013 -925 2015
rect 896 2012 898 2014
rect 896 1992 898 1994
rect 896 1972 898 1974
rect -891 1922 -889 1924
rect -891 1812 -889 1814
rect 896 1812 898 1814
rect 896 1792 898 1794
rect 829 1780 831 1782
rect 834 1780 836 1782
rect 839 1780 841 1782
rect 829 1775 831 1777
rect 834 1775 836 1777
rect 839 1775 841 1777
rect 829 1770 831 1772
rect 834 1770 836 1772
rect 839 1770 841 1772
rect 829 1765 831 1767
rect 834 1765 836 1767
rect 839 1765 841 1767
rect 829 1760 831 1762
rect 834 1760 836 1762
rect 839 1760 841 1762
rect 829 1755 831 1757
rect 834 1755 836 1757
rect 839 1755 841 1757
rect 829 1750 831 1752
rect 834 1750 836 1752
rect 839 1750 841 1752
rect 829 1745 831 1747
rect 834 1745 836 1747
rect 839 1745 841 1747
rect 829 1740 831 1742
rect 834 1740 836 1742
rect 839 1740 841 1742
rect 829 1735 831 1737
rect 834 1735 836 1737
rect 839 1735 841 1737
rect 829 1730 831 1732
rect 834 1730 836 1732
rect 839 1730 841 1732
rect 829 1725 831 1727
rect 834 1725 836 1727
rect 839 1725 841 1727
rect 829 1720 831 1722
rect 834 1720 836 1722
rect 839 1720 841 1722
rect 829 1715 831 1717
rect 834 1715 836 1717
rect 839 1715 841 1717
rect 829 1710 831 1712
rect 834 1710 836 1712
rect 839 1710 841 1712
rect -891 1692 -889 1694
rect -891 1492 -889 1494
rect -890 1292 -888 1294
rect -891 1242 -889 1244
rect -1492 -688 -1490 -686
rect -1490 -988 -1488 -986
rect -1492 -1288 -1490 -1286
rect 112 -1376 114 -1374
rect 23 -1384 25 -1382
rect -1388 -1391 -1386 -1389
rect -1088 -1390 -1086 -1388
rect 412 -1389 414 -1387
rect -788 -1392 -786 -1390
rect 712 -1392 714 -1390
rect 1012 -1391 1014 -1389
rect 1312 -1392 1314 -1390
rect 2211 -1391 2213 -1389
rect 1911 -1393 1913 -1391
<< metal3 >>
rect -1489 3358 -1324 3364
rect -1330 3195 -1324 3358
rect -1242 3225 -1233 3385
rect -942 3241 -933 3386
rect -642 3257 -633 3386
rect -342 3272 -333 3386
rect -42 3288 -33 3386
rect 258 3304 267 3389
rect 858 3320 867 3386
rect 1158 3320 1167 3386
rect 1456 3343 1466 3385
rect 858 3312 936 3320
rect 978 3312 1167 3320
rect 1365 3333 1468 3343
rect 258 3296 924 3304
rect -42 3280 948 3288
rect -343 3264 996 3272
rect -642 3249 95 3257
rect -942 3233 -17 3241
rect -226 3232 -17 3233
rect -1242 3217 -345 3225
rect -1330 3185 -886 3195
rect -1445 3056 -898 3066
rect -1445 2756 -910 2766
rect -1445 2456 -934 2465
rect -955 2016 -949 2017
rect -1439 2011 -946 2016
rect -1439 1633 -1433 2011
rect -940 1946 -934 2456
rect -916 2036 -910 2756
rect -904 2226 -898 3056
rect -892 2556 -886 3185
rect -351 2751 -345 3217
rect -22 2892 -17 3232
rect -23 2751 -17 2892
rect 89 2751 95 3249
rect -892 2551 -866 2556
rect -904 2221 -866 2226
rect 894 2077 900 2864
rect 877 2071 900 2077
rect -886 2056 -880 2057
rect 889 2056 895 2057
rect -892 2051 -867 2056
rect 878 2051 900 2056
rect -916 2031 -866 2036
rect 877 2031 900 2037
rect -925 2016 -919 2017
rect 889 2016 895 2017
rect -928 2011 -866 2016
rect 878 2011 900 2016
rect 889 1996 895 1997
rect 878 1991 900 1996
rect 889 1976 895 1977
rect 878 1971 900 1976
rect 918 1957 924 3252
rect 877 1951 924 1957
rect -940 1941 -866 1946
rect 930 1937 936 3252
rect 877 1931 936 1937
rect -892 1921 -866 1926
rect -889 1920 -883 1921
rect 942 1917 948 3252
rect 990 3251 996 3264
rect 878 1911 948 1917
rect 954 3207 1327 3215
rect 954 1897 960 3207
rect 1365 3199 1375 3333
rect 1758 3215 1766 3386
rect 1396 3207 1766 3215
rect 2055 3385 2060 3387
rect 878 1891 960 1897
rect 966 3191 1375 3199
rect 966 1877 972 3191
rect 878 1871 972 1877
rect 978 1857 984 3119
rect 882 1851 984 1857
rect 990 1837 996 3119
rect 2055 3065 2064 3385
rect 1028 3056 2064 3065
rect 1028 2864 1034 3056
rect 1007 2857 1034 2864
rect -1424 1831 -866 1836
rect 882 1831 996 1837
rect -1424 1565 -1418 1831
rect 889 1816 895 1817
rect -892 1811 -866 1816
rect 878 1811 900 1816
rect -889 1810 -883 1811
rect 889 1796 895 1797
rect 878 1791 900 1796
rect -892 1691 -866 1696
rect -889 1690 -883 1691
rect -1445 1556 -1418 1565
rect -1402 1631 -866 1636
rect -1402 1265 -1390 1631
rect -1445 1256 -1390 1265
rect -1370 1541 -866 1546
rect -1370 965 -1361 1541
rect -892 1491 -866 1496
rect -889 1490 -883 1491
rect -1445 956 -1361 965
rect -1334 1341 -866 1346
rect -1334 665 -1324 1341
rect -1445 656 -1324 665
rect -1299 1321 -866 1326
rect -1299 542 -1289 1321
rect -892 1291 -866 1296
rect -888 1290 -882 1291
rect -892 1241 -866 1246
rect -889 1240 -883 1241
rect -1299 530 -1233 542
rect -1242 -157 -1233 530
rect -1490 -166 -1233 -157
rect -1242 -171 -1233 -166
<< gv2 >>
rect -939 3382 -937 3384
rect -639 3382 -637 3384
rect -338 3382 -336 3384
rect -38 3382 -36 3384
rect 262 3383 264 3385
rect 862 3382 864 3384
rect 1161 3382 1163 3384
rect -1239 3380 -1237 3382
rect 1460 3381 1462 3383
rect 1761 3382 1763 3384
rect 2058 3381 2060 3383
rect -1487 3360 -1485 3362
rect 932 3315 934 3317
rect 980 3315 982 3317
rect 920 3299 922 3301
rect 944 3283 946 3285
rect 992 3258 994 3260
rect 992 3253 994 3255
rect 932 3248 934 3250
rect 944 3248 946 3250
rect 920 3246 922 3248
rect 932 3243 934 3245
rect 944 3243 946 3245
rect 920 3241 922 3243
rect 932 3238 934 3240
rect 944 3238 946 3240
rect 1317 3210 1319 3212
rect 1322 3210 1324 3212
rect 1398 3210 1400 3212
rect 1403 3210 1405 3212
rect 980 3110 982 3112
rect 992 3110 994 3112
rect -1441 3059 -1439 3061
rect 896 2859 898 2861
rect 1011 2859 1013 2861
rect -1440 2760 -1438 2762
rect -349 2753 -347 2755
rect -21 2753 -19 2755
rect 91 2753 93 2755
rect -1441 2459 -1439 2461
rect -884 2053 -882 2055
rect 891 2053 893 2055
rect 891 2033 893 2035
rect -953 2013 -951 2015
rect -923 2013 -921 2015
rect 891 2013 893 2015
rect 891 1993 893 1995
rect 891 1973 893 1975
rect -887 1922 -885 1924
rect -887 1812 -885 1814
rect 891 1813 893 1815
rect 891 1793 893 1795
rect -887 1692 -885 1694
rect -1437 1636 -1435 1638
rect -1440 1559 -1438 1561
rect -887 1492 -885 1494
rect -886 1292 -884 1294
rect -1441 1259 -1439 1261
rect -887 1242 -885 1244
rect -1440 959 -1438 961
rect -1441 659 -1439 661
rect -1487 -163 -1485 -161
use PadFC  16_0
timestamp 1683038052
transform 1 0 -2500 0 1 3400
box 330 -3 1003 670
use PadBiDir  17_0
timestamp 1683038052
transform 1 0 -1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_1
timestamp 1683038052
transform 1 0 -1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_2
timestamp 1683038052
transform 1 0 -900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_3
timestamp 1683038052
transform 1 0 -600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_4
timestamp 1683038052
transform 1 0 -300 0 1 3400
box -36 -19 303 1000
use PadVdd  18_0
timestamp 1683038052
transform 1 0 300 0 1 3400
box -3 -12 303 1000
use PadBiDir  17_5
timestamp 1683038052
transform 1 0 0 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_6
timestamp 1683038052
transform 1 0 600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_7
timestamp 1683038052
transform 1 0 900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_8
timestamp 1683038052
transform 1 0 1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_0
timestamp 1683038052
transform 1 0 1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_1
timestamp 1683038052
transform 1 0 1800 0 1 3400
box -36 -19 303 1000
use PadVdd  PadVdd_0
timestamp 1683038052
transform 1 0 2400 0 1 3400
box -3 -12 303 1000
use PadBiDir  PadBiDir_2
timestamp 1683038052
transform 1 0 2100 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_3
timestamp 1683038052
transform 1 0 2700 0 1 3400
box -36 -19 303 1000
use PadFC  16_1
timestamp 1683038052
transform 0 1 3300 -1 0 4400
box 330 -3 1003 670
use PadBiDir  PadBiDir_4
timestamp 1683038052
transform 1 0 3000 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_9
timestamp 1683038052
transform 0 -1 -1500 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_10
timestamp 1683038052
transform 0 -1 -1500 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_17
timestamp 1683038052
transform 0 1 3300 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_18
timestamp 1683038052
transform 0 1 3300 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_11
timestamp 1683038052
transform 0 -1 -1500 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_12
timestamp 1683038052
transform 0 -1 -1500 1 0 2200
box -36 -19 303 1000
use PadGnd  19_0
timestamp 1683038052
transform 0 -1 -1500 -1 0 2200
box -3 -11 303 1000
use PadBiDir  17_13
timestamp 1683038052
transform 0 -1 -1500 -1 0 1900
box -36 -19 303 1000
use PadBiDir  PadBiDir_14
timestamp 1683038052
transform 0 -1 -1500 1 0 1300
box -36 -19 303 1000
use CORDIC_TOP  CORDIC_TOP_0
timestamp 1683038052
transform 1 0 -880 0 1 1019
box 0 13 1767 1740
use PadBiDir  17_19
timestamp 1683038052
transform 0 1 3300 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_20
timestamp 1683038052
transform 0 1 3300 1 0 2200
box -36 -19 303 1000
use PadBiDir  17_21
timestamp 1683038052
transform 0 1 3300 1 0 1900
box -36 -19 303 1000
use PadGnd  19_1
timestamp 1683038052
transform 0 1 3300 -1 0 1900
box -3 -11 303 1000
use PadBiDir  PadBiDir_19
timestamp 1683038052
transform 0 1 3300 1 0 1300
box -36 -19 303 1000
use PadBiDir  PadBiDir_13
timestamp 1683038052
transform 0 -1 -1500 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_12
timestamp 1683038052
transform 0 -1 -1500 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_11
timestamp 1683038052
transform 0 -1 -1500 1 0 400
box -36 -19 303 1000
use PadBiDir  PadBiDir_18
timestamp 1683038052
transform 0 1 3300 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_17
timestamp 1683038052
transform 0 1 3300 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_16
timestamp 1683038052
transform 0 1 3300 1 0 400
box -36 -19 303 1000
use PadGnd  PadGnd_0
timestamp 1683038052
transform 0 -1 -1500 -1 0 400
box -3 -11 303 1000
use PadBiDir  PadBiDir_15
timestamp 1683038052
transform 0 1 3300 1 0 100
box -36 -19 303 1000
use PadBiDir  PadBiDir_10
timestamp 1683038052
transform 0 -1 -1500 -1 0 100
box -36 -19 303 1000
use PadBiDir  17_14
timestamp 1683038052
transform 0 -1 -1500 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_15
timestamp 1683038052
transform 0 -1 -1500 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_16
timestamp 1683038052
transform 0 -1 -1500 1 0 -1100
box -36 -19 303 1000
use PadGnd  PadGnd_1
timestamp 1683038052
transform 0 1 3300 -1 0 100
box -3 -11 303 1000
use PadBiDir  17_22
timestamp 1683038052
transform 0 1 3300 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_23
timestamp 1683038052
transform 0 1 3300 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_24
timestamp 1683038052
transform 0 1 3300 1 0 -1100
box -36 -19 303 1000
use PadBiDir  17_25
timestamp 1683038052
transform 0 -1 -1500 1 0 -1400
box -36 -19 303 1000
use PadFC  16_2
timestamp 1683038052
transform 0 -1 -1500 1 0 -2400
box 330 -3 1003 670
use PadBiDir  17_26
timestamp 1683038052
transform 1 0 -1500 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_27
timestamp 1683038052
transform 1 0 -1200 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_28
timestamp 1683038052
transform 1 0 -900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_29
timestamp 1683038052
transform 1 0 -600 0 -1 -1400
box -36 -19 303 1000
use PadVdd  18_1
timestamp 1683038052
transform 1 0 -300 0 -1 -1400
box -3 -12 303 1000
use PadBiDir  17_30
timestamp 1683038052
transform 1 0 0 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_31
timestamp 1683038052
transform 1 0 300 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_32
timestamp 1683038052
transform 1 0 600 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_33
timestamp 1683038052
transform 1 0 900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_35
timestamp 1683038052
transform 1 0 1200 0 -1 -1400
box -36 -19 303 1000
use PadVdd  PadVdd_1
timestamp 1683038052
transform 1 0 1500 0 -1 -1400
box -3 -12 303 1000
use PadBiDir  PadBiDir_5
timestamp 1683038052
transform 1 0 1800 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_6
timestamp 1683038052
transform 1 0 2100 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_7
timestamp 1683038052
transform 1 0 2400 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_8
timestamp 1683038052
transform 1 0 2700 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_34
timestamp 1683038052
transform 0 1 3300 1 0 -1400
box -36 -19 303 1000
use PadFC  16_3
timestamp 1683038052
transform -1 0 4300 0 -1 -1400
box 330 -3 1003 670
use PadBiDir  PadBiDir_9
timestamp 1683038052
transform 1 0 3000 0 -1 -1400
box -36 -19 303 1000
<< labels >>
rlabel metal1 -1352 4113 -1352 4113 4 p_clkb
rlabel metal1 -1052 4111 -1052 4111 4 p_clka
rlabel metal1 -751 4115 -751 4115 4 p_in_port0_0
rlabel metal1 -455 4108 -455 4108 4 p_in_port0_1
rlabel metal1 -138 4113 -138 4113 4 p_in_port0_2
rlabel metal1 149 4102 149 4102 6 p_in_port0_3
rlabel metal1 739 4111 739 4111 6 p_in_port0_4
rlabel metal1 1046 4120 1046 4120 6 p_in_port0_5
rlabel metal1 1334 4104 1334 4104 6 p_in_port0_6
rlabel metal1 1652 4117 1652 4117 6 p_in_port0_7
rlabel metal1 1940 4100 1940 4100 6 p_cordic_mode
rlabel metal1 -2208 2655 -2208 2655 4 p_in_port1_7
rlabel metal1 -2210 2357 -2210 2357 4 p_in_port1_6
rlabel metal1 -2217 1746 -2217 1746 4 p_in_port1_5
rlabel metal1 -2215 1447 -2215 1447 4 p_in_port1_4
rlabel metal1 -2208 1156 -2208 1156 4 p_in_port1_3
rlabel metal1 -2204 843 -2204 843 4 p_in_port1_2
rlabel metal1 -2208 550 -2208 550 4 p_in_port1_1
rlabel metal1 -2217 -41 -2217 -41 2 p_in_port1_0
rlabel metal1 -2204 -354 -2204 -354 2 p_out_port1_5
rlabel metal1 -2208 -656 -2208 -656 2 p_out_port1_6
rlabel metal1 -2204 -945 -2204 -945 2 p_out_port1_4
rlabel metal1 -1047 -2110 -1047 -2110 2 p_out_port1_3
rlabel metal1 -750 -2106 -750 -2106 2 p_out_port1_2
rlabel metal1 -455 -2108 -455 -2108 2 p_out_port1_1
rlabel metal1 138 -2103 138 -2103 8 p_out_port1_0
rlabel metal1 456 -2106 456 -2106 8 p_out_port0_6
rlabel metal1 751 -2115 751 -2115 8 p_out_port0_7
rlabel metal1 1055 -2106 1055 -2106 8 p_out_port0_5
rlabel metal1 1364 -2103 1364 -2103 8 p_out_port0_4
rlabel metal1 1939 -2108 1939 -2108 8 p_out_port0_2
rlabel metal1 2250 -2110 2250 -2110 8 p_out_port0_3
rlabel metal1 2541 -2106 2541 -2106 8 p_out_port0_1
rlabel metal1 4002 3255 4002 3255 6 p_done
rlabel metal1 4007 2957 4007 2957 6 p_out_port1_7
rlabel metal1 4016 2663 4016 2663 6 p_out_port0_0
rlabel metal1 -2210 3254 -2210 3254 4 p_reset
rlabel metal1 -2213 2945 -2213 2945 4 p_start
rlabel metal2 909 1974 909 1974 6 out_port0_5
rlabel metal1 446 4106 446 4106 6 Vdd
rlabel metal1 -2210 2051 -2210 2051 4 GND
rlabel metal3 903 1833 903 1833 6 in_port0_1
rlabel metal3 903 1854 903 1854 6 in_port0_5
rlabel metal3 902 1873 902 1873 6 in_port0_6
rlabel metal3 900 1894 900 1894 6 in_port0_7
rlabel metal3 899 1912 899 1912 6 in_port0_2
rlabel metal3 899 1933 899 1933 6 in_port0_4
rlabel metal3 899 1954 899 1954 6 in_port0_3
rlabel metal3 896 2074 896 2074 6 cordic_mode
rlabel metal3 -348 2753 -348 2753 4 clkb
rlabel metal3 92 2754 92 2754 6 in_port0_0
rlabel metal3 -20 2753 -20 2753 4 clka
rlabel metal3 -873 2554 -873 2554 4 reset
rlabel metal3 -872 2223 -872 2223 4 start
rlabel metal3 -870 2033 -870 2033 4 in_port1_7
rlabel metal3 -870 2014 -870 2014 4 in_port1_5
rlabel metal3 -870 1943 -870 1943 4 in_port1_6
rlabel metal3 -870 1833 -870 1833 4 in_port1_4
rlabel metal3 -869 1632 -869 1632 4 in_port1_3
rlabel metal3 -869 1543 -869 1543 4 in_port1_2
rlabel metal3 -869 1343 -869 1343 4 in_port1_1
rlabel metal3 -868 1324 -868 1324 4 in_port1_0
<< end >>
