magic
tech scmos
timestamp 1681696376
<< nwell >>
rect -5 48 28 105
<< ntransistor >>
rect 7 6 9 16
rect 15 6 17 26
<< ptransistor >>
rect 7 74 9 94
rect 15 54 17 94
<< ndiffusion >>
rect 10 25 15 26
rect 2 15 7 16
rect 6 6 7 15
rect 9 6 10 16
rect 14 6 15 25
rect 17 25 22 26
rect 17 6 18 25
<< pdiffusion >>
rect 2 93 7 94
rect 6 74 7 93
rect 9 74 10 94
rect 14 60 15 94
rect 10 54 15 60
rect 17 93 22 94
rect 17 54 18 93
<< ndcontact >>
rect 2 6 6 15
rect 10 6 14 25
rect 18 6 22 25
<< pdcontact >>
rect 2 74 6 93
rect 10 60 14 94
rect 18 54 22 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 7 57 9 74
rect 6 55 9 57
rect 6 41 8 55
rect 15 51 17 54
rect 16 47 17 51
rect 6 39 9 41
rect 7 16 9 39
rect 15 26 17 47
rect 7 4 9 6
rect 15 4 17 6
<< polycontact >>
rect 2 39 6 43
rect 12 47 16 51
<< metal1 >>
rect -2 102 26 103
rect 2 98 14 102
rect 18 98 26 102
rect -2 97 26 98
rect 10 94 14 97
rect 2 93 6 94
rect 2 57 6 74
rect 18 93 22 94
rect 2 54 13 57
rect 10 51 13 54
rect 10 47 12 51
rect 2 43 6 47
rect 10 32 13 47
rect 19 43 22 54
rect 2 29 13 32
rect 2 15 6 29
rect 10 25 14 26
rect 18 25 22 43
rect 10 3 14 6
rect -2 2 26 3
rect 2 -2 14 2
rect 18 -2 26 2
rect -2 -3 26 -2
<< m1p >>
rect 2 43 6 47
rect 18 33 22 37
<< labels >>
rlabel metal1 4 100 4 100 4 vdd
rlabel metal1 4 0 4 0 4 gnd
rlabel metal1 4 45 4 45 4 A
rlabel metal1 20 35 20 35 4 Y
<< end >>
