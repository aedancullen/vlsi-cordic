magic
tech scmos
timestamp 1681696376
<< m2contact >>
rect -2 -2 2 2
<< end >>
