magic
tech scmos
timestamp 1683038052
<< nwell >>
rect -5 48 53 105
rect 6 44 33 48
<< ntransistor >>
rect 7 10 9 20
rect 15 10 17 30
rect 20 10 22 30
rect 28 10 30 30
rect 33 10 35 30
<< ptransistor >>
rect 7 70 9 90
rect 15 50 17 90
rect 20 50 22 90
rect 28 54 30 94
rect 33 54 35 94
<< ndiffusion >>
rect 12 28 15 30
rect 10 20 15 28
rect 2 10 7 20
rect 9 10 15 20
rect 17 10 20 30
rect 22 10 28 30
rect 30 10 33 30
rect 35 10 40 30
<< pdiffusion >>
rect 23 90 28 94
rect 2 70 7 90
rect 9 70 15 90
rect 10 56 15 70
rect 12 50 15 56
rect 17 50 20 90
rect 22 54 28 90
rect 30 54 33 94
rect 35 54 40 94
rect 22 50 25 54
<< psubstratepdiff >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
<< nsubstratendiff >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
<< polysilicon >>
rect 7 95 22 97
rect 7 90 9 95
rect 15 90 17 92
rect 20 90 22 95
rect 28 94 30 96
rect 33 94 35 96
rect 7 69 9 70
rect 4 67 9 69
rect 4 43 6 67
rect 15 49 17 50
rect 12 47 17 49
rect 20 48 22 50
rect 12 43 14 47
rect 2 39 6 43
rect 10 39 14 43
rect 28 40 30 54
rect 33 53 35 54
rect 33 51 36 53
rect 4 23 6 39
rect 11 33 13 39
rect 21 38 30 40
rect 34 47 38 51
rect 21 36 25 38
rect 20 34 24 36
rect 11 31 17 33
rect 15 30 17 31
rect 20 30 22 34
rect 34 33 36 47
rect 28 30 30 32
rect 33 31 36 33
rect 33 30 35 31
rect 4 21 9 23
rect 7 20 9 21
rect 7 5 9 10
rect 15 8 17 10
rect 20 8 22 10
rect 28 5 30 10
rect 33 8 35 10
rect 7 3 30 5
<< genericcontact >>
rect -1 99 1 101
rect 15 99 17 101
rect 31 99 33 101
rect 24 89 26 91
rect 37 90 39 92
rect 3 86 5 88
rect 11 87 13 89
rect 24 84 26 86
rect 37 85 39 87
rect 3 81 5 83
rect 11 82 13 84
rect 24 79 26 81
rect 37 80 39 82
rect 3 76 5 78
rect 11 77 13 79
rect 24 74 26 76
rect 37 75 39 77
rect 3 71 5 73
rect 11 72 13 74
rect 24 69 26 71
rect 37 70 39 72
rect 11 67 13 69
rect 24 64 26 66
rect 37 65 39 67
rect 11 62 13 64
rect 24 59 26 61
rect 37 60 39 62
rect 11 57 13 59
rect 37 55 39 57
rect 35 48 37 50
rect 3 40 5 42
rect 11 40 13 42
rect 22 37 24 39
rect 37 26 39 28
rect 11 23 13 25
rect 24 23 26 25
rect 37 21 39 23
rect 11 18 13 20
rect 24 18 26 20
rect 3 16 5 18
rect 37 16 39 18
rect 11 13 13 15
rect 24 13 26 15
rect 3 11 5 13
rect 37 11 39 13
rect -1 -1 1 1
rect 15 -1 17 1
rect 31 -1 33 1
<< metal1 >>
rect -2 97 50 103
rect 2 70 6 90
rect 2 53 5 70
rect 10 56 14 97
rect 23 59 27 94
rect 23 56 31 59
rect 2 50 21 53
rect 2 39 6 47
rect 10 39 14 47
rect 18 40 21 50
rect 18 36 25 40
rect 28 37 31 56
rect 36 54 40 97
rect 34 43 38 51
rect 18 34 23 36
rect 2 31 23 34
rect 28 33 38 37
rect 2 20 5 31
rect 28 30 31 33
rect 27 28 31 30
rect 2 10 6 20
rect 10 3 14 28
rect 23 25 31 28
rect 23 10 27 25
rect 36 3 40 30
rect -2 -3 50 3
<< m1p >>
rect 2 43 6 47
rect 10 43 14 47
rect 34 43 38 47
rect 34 33 38 37
<< labels >>
rlabel metal1 4 45 4 45 6 S
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 36 35 36 35 6 Y
rlabel metal1 36 45 36 45 6 A
rlabel metal1 12 45 12 45 6 B
<< end >>
